--
-- FB_top.vhd
-- Author : David Humphrey (dave.humphrey@csiro.au)
-- Description
--  Top level for the correlator filterbanks. Includes :
--   - Correlator filterbank - 4096 point FFT, 12 tap FIR filter, 4 streams simultaneously.
--   - Fine delay
--   - MACE interface, which is just to allow reading/writing of the filter taps in the filterbanks.
--     *** WARNING *** MACE slave is manually written. MACE slave module is NOT auto-generated by ARGS. 
--     Changing the yaml file will not change the actual registers.
--     This is to allow the memories to reside in the filters, rather than being pulled out and put into 
--     ARGs. 
--
----------------------------------------------------------------------------------------------------------
library IEEE, axi4_lib, common_lib, filterbanks_lib, dsp_top_lib;

use dsp_top_lib.dsp_top_pkg.all;
use common_lib.common_pkg.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use axi4_lib.axi4_lite_pkg.ALL;
use axi4_lib.axi4_full_pkg.ALL;
Library xpm;
use xpm.vcomponents.all;
USE filterbanks_lib.cor_filterbanks_filterbanks_reg_pkg.ALL;

entity FB_Top_correlator_dummy is
    port(
        i_data_rst  : in std_logic;
        -- AXI slave interface, 64k word block of space with the fir filter coefficients.
        i_axi_clk  : in std_logic;
        i_axi_rst  : in std_logic;
        i_axi_mosi  : in  t_axi4_lite_mosi;
        o_axi_miso  : out t_axi4_lite_miso;
        -- Configuration (on i_data_clk)
        i_fineDelayDisable : in std_logic;
        -----------------------------------------
        -- data input, common valid signal, expects packets of 64 samples. 
        -- Requires at least 2 clocks idle time between packets.
        i_SOF    : in std_logic; 
        i_data0  : in t_slv_16_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        i_data1  : in t_slv_16_arr(1 downto 0);
        i_meta01 : in t_CT1_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(31:0), virtualChannel(15:0), .valid
        i_data2  : in t_slv_16_arr(1 downto 0);
        i_data3  : in t_slv_16_arr(1 downto 0);
        i_meta23 : in t_CT1_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(31:0), virtualChannel(15:0), .valid
        i_data4  : in t_slv_16_arr(1 downto 0);
        i_data5  : in t_slv_16_arr(1 downto 0);
        i_meta45 : in t_CT1_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(31:0), virtualChannel(15:0), .valid
        i_data6  : in t_slv_16_arr(1 downto 0);
        i_data7  : in t_slv_16_arr(1 downto 0);
        i_meta67 : in t_CT1_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(31:0), virtualChannel(15:0), .valid
        --
        i_lastChannel : in std_logic;
        i_demap_table_select : in std_logic;
        --
        i_DataValid : in std_logic;
        -- Correlator filterbank data output
        o_integration    : out std_logic_vector(31 downto 0); -- integration in units of 849ms since epoch.
        o_ctFrame        : out std_logic_vector(1 downto 0); -- corner turn frame, 0, 1 or 2, units of 283ms relative to integration.
        o_virtualChannel : out t_slv_16_arr(3 downto 0); -- 3 virtual channels, one for each of the PST data streams.
        o_bad_poly       : out std_logic;
        --
        o_lastChannel    : out std_logic;  -- Last of the group of 4 channels
        o_demap_table_select : out std_logic;
        --
        o_HeaderValid : out std_logic_vector(3 downto 0);
        o_Data        : out t_ctc_output_payload_arr(3 downto 0);
        o_DataValid   : out std_logic;
        -- i_SOF delayed by 16384 clocks;
        -- i_sof occurs at the start of each new block of 4 virtual channels.
        -- Delay of 16384 is enough to ensure that o_sof falls in the gap
        -- between data packets at the filterbank output that occurs due to the filterbank preload.
        o_sof : out std_logic;
        -- Correlator filterbank output as packets
        -- Each output packet contains all the data for:
        --  - Single time step
        --  - Single polarisation
        --  - single coarse channel
        -- This is 3456 * 2 (re+im) bytes, plus 16 bytes of header.
        -- The data is transferred in bursts of 433 clocks.
        o_packetData : out std_logic_vector(127 downto 0);
        o_packetValid : out std_logic;
        i_packetReady : in std_logic
    );

    -- prevent optimisation across module boundaries.
    attribute keep_hierarchy : string;
    attribute keep_hierarchy of FB_Top_correlator_dummy : entity is "yes";
    
end FB_Top_correlator_dummy;

architecture Behavioral of FB_Top_correlator_dummy is
    
    signal FDdata  : t_ctc_output_payload_arr(3 downto 0);
    
    signal firtap_addr : std_logic_vector(15 downto 0);
    --signal firtap_clk : std_logic;
    signal cor_we : std_logic;
    signal corFirRd_data : std_logic_vector(17 downto 0);
    signal firtap_wr_data : std_logic_vector(17 downto 0);
    
    signal CorDin0, CorDin1, CorDin2, CorDin3 : t_slv_8_arr(1 downto 0);
    signal CorrelatorMetaIn, CorrelatorMetaOut : std_logic_vector(619 downto 0);
    signal CorDout0, CorDout1, CorDout2, CorDout3 : t_slv_16_arr(1 downto 0);
    signal CorValidOut, CorValidOutDel : std_logic;
    
    signal data0, data1, data2, data3, data4, data5, data6, data7 : t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.  
    
    signal FDcorDataValid : std_logic_vector(3 downto 0);
    
    signal corFBHeader : t_CT1_META_out_arr(3 downto 0);
    signal corDout_arr : t_FB_output_payload_a(3 downto 0);
    
    signal FDHeader : t_CT1_META_out_arr(3 downto 0);
    signal DataValid : std_logic;
    
    signal corFBDout0, corFBDout1, corFBDout2, corFBDout3, corFBDout4, corFBDout5, corFBDout6, corFBDout7, corFBDout8 : t_slv_16_arr(1 downto 0);
    signal corMetaOut : std_logic_vector(619 downto 0);
    
    signal corFBHeaderValid : std_logic;
    
    signal captureCount : std_logic_vector(3 downto 0);
    signal FDcorDataValidDel1 : std_logic;
    signal captureData : t_slv_256_arr(7 downto 0);
    
    signal triggerRdLow128bits : std_logic_vector(6 downto 0) := "0000000";
    signal triggerRdHigh128bits : std_logic_vector(6 downto 0) := "0000000";
    signal copyToUramCount : std_logic_Vector(2 downto 0);
    signal copyToUramValidLow, copyToUramValidHigh, copyToUramValidLowDel1, copyToUramValidHighDel1 : std_logic := '0';
    signal bufWrAddrDoubleBufferSelect : std_logic := '0';
    signal bufWrAddrBuffer, bufWrAddrBufferAdv : std_logic_vector(2 downto 0);
    signal bufWrAddrWord : std_logic_vector(8 downto 0);
    signal bufRdAddrDoubleBufferSelect : std_logic := '0';
    signal bufRdAddrBuffer, bufRdAddrBufferDel1, bufRdAddrBufferDel2, bufRdAddrBufferDel3 : std_logic_vector(2 downto 0);
    signal bufRdAddrWord : std_logic_vector(8 downto 0);
    signal bufWE : std_logic_vector(0 downto 0);
    type sendTo100GE_fsm_t is (start, checkEnable, checkEnableWait0, checkEnableWait1, checkEnableWait2, checkEnableWait3, waitReady, sendHeader, sendData, nextBuffer, done);
    signal sendTo100GE_fsm : sendTo100GE_fsm_t := done;
    signal sendTo100GE_fsm_del1, sendTo100GE_fsm_del2, sendTo100GE_fsm_del3 : sendTo100GE_fsm_t := done;

    signal bufWrData, bufDout : std_logic_vector(127 downto 0);
    signal triggerSendTo100GE : std_logic;
    signal vc_hold, vc_out : t_slv_16_arr(3 downto 0);
    signal framecount_hold, framecount_out : std_logic_vector(31 downto 0);
    signal bufWrAddr, bufRdAddr : std_logic_vector(12 downto 0);
    signal config_ro : t_config_ro;
    signal output_disable_i : t_config_output_disable_ram_in;
    signal output_disable_o : t_config_output_disable_ram_out;
    signal tx_packet_count, tx_packet_count_ct : std_logic_vector(31 downto 0) := x"00000000";
    signal packetValidDel1, packetValid, FDcorDataValidDel : std_logic;
    signal output_disabled : std_logic;
    signal output_disable_addr : std_logic_vector(9 downto 0);
    signal reg_reset_del1, reg_reset : std_logic;
    signal config_rw : t_config_rw;
    signal HeaderValid : std_logic_vector(3 downto 0);
    signal sof_out, sof_del1 : std_logic := '0';
    signal sof_out_count : std_logic_vector(13 downto 0) := (others => '0');
    
    signal FD_datavalid, FD_headerValid : std_logic_vector(18 downto 0);
    signal FD_finecount : std_logic_vector(15 downto 0);
    signal FD_virtualChannel0, FD_virtualChannel1, FD_virtualChannel2, FD_virtualChannel3 : t_slv_16_arr(18 downto 0);
    signal FD_integration : t_slv_32_arr(18 downto 0);
    signal FD_ctFrame : t_slv_2_arr(18 downto 0);
    signal FD_bad_poly, FD_lastChannel, FD_demap_table_select : std_logic_vector(18 downto 0);
    
begin
    
    -----------------------------------------------------------------------------------
    -- correlator Filterbank
    process(i_axi_clk)
    begin
        if rising_edge(i_axi_clk) then
            CorrelatorMetaIn(31 downto 0)               <= i_meta01.HDeltaP;
            CorrelatorMetaIn(63 downto 32)              <= i_meta01.VDeltaP;
            CorrelatorMetaIn(95 downto 64)              <= i_meta01.HOffsetP;
            CorrelatorMetaIn(127 downto 96)             <= i_meta01.VOffsetP;
            CorrelatorMetaIn(143 downto 128)            <= i_meta01.virtualChannel;
            CorrelatorMetaIn(144)                       <= i_meta01.valid; -- note that .valid is just a qualifier for the meta data. The meta data is only valid if both this and i_datavalid are high.
            
            CorrelatorMetaIn(31+145 downto 0+145)       <= i_meta23.HDeltaP;
            CorrelatorMetaIn(63+145 downto 32+145)      <= i_meta23.VDeltaP;
            CorrelatorMetaIn(95+145 downto 64+145)      <= i_meta23.HOffsetP;
            CorrelatorMetaIn(127+145 downto 96+145)     <= i_meta23.VOffsetP;
            CorrelatorMetaIn(143+145 downto 128+145)    <= i_meta23.virtualChannel;
            CorrelatorMetaIn(144+145)                   <= i_meta23.valid;
            
            CorrelatorMetaIn(31+290 downto 0+290)       <= i_meta45.HDeltaP;
            CorrelatorMetaIn(63+290 downto 32+290)      <= i_meta45.VDeltaP;
            CorrelatorMetaIn(95+290 downto 64+290)      <= i_meta45.HOffsetP;
            CorrelatorMetaIn(127+290 downto 96+290)     <= i_meta45.VOffsetP;
            CorrelatorMetaIn(143+290 downto 128+290)    <= i_meta45.virtualChannel;
            CorrelatorMetaIn(144+290)                   <= i_meta45.valid;

            CorrelatorMetaIn(31+435 downto 0+435)       <= i_meta67.HDeltaP;
            CorrelatorMetaIn(63+435 downto 32+435)      <= i_meta67.VDeltaP;
            CorrelatorMetaIn(95+435 downto 64+435)      <= i_meta67.HOffsetP;
            CorrelatorMetaIn(127+435 downto 96+435)     <= i_meta67.VOffsetP;
            CorrelatorMetaIn(143+435 downto 128+435)    <= i_meta67.virtualChannel;
            CorrelatorMetaIn(144+435)                   <= i_meta67.valid;
            
            CorrelatorMetaIn(31+580 downto 0+580)       <= i_meta01.integration;  -- framecount is the same for all input headers. Total of 32+4*81 = 356 header bits.
            CorrelatorMetaIn(33+580 downto 32+580)      <= i_meta01.ctFrame;
            
            CorrelatorMetaIn(614) <= i_meta01.bad_poly;
            CorrelatorMetaIn(615) <= i_meta23.bad_poly;
            CorrelatorMetaIn(616) <= i_meta45.bad_poly;
            CorrelatorMetaIn(617) <= i_meta67.bad_poly;
            CorrelatorMetaIn(618) <= i_lastChannel;
            CorrelatorMetaIn(619) <= i_demap_table_select;
            DataValid <= i_DataValid;
            
            -- Generate o_sof from i_sof, taking into account the latency of the filterbank processing.
            sof_del1 <= i_sof;
            if i_sof = '1' and sof_del1 = '0' then
                sof_out_count <= (others => '1'); -- 16383
            elsif (unsigned(sof_out_count) /= 0) then
                sof_out_count <= std_logic_vector(unsigned(sof_out_count) - 1);
            end if;
            if (unsigned(sof_out_count) = 1) then
                sof_out <= '1';
            else
                sof_out <= '0';
            end if;
            o_sof <= sof_out;
        end if;
    end process;
    
    
--    corfbi : entity filterbanks_lib.correlatorFBTop25
--    generic map(
--        METABITS => 361,    -- Width in bits of the meta_i and meta_o ports.
--        FRAMESTODROP => 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
--    ) port map (
--        -- processing clock
--        clk     => i_axi_clk,
--        rst     => i_SOF,
--        -- Data input, common valid signal, expects packets of 64 samples. 
--        -- Requires at least 2 clocks idle time between packets.
--        -- Due to oversampling, also requires on average 86 clocks between packets - specifically, no more than 3 packets in 258 clocks. 
--        data0_i => data0, -- in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
--        data1_i => data1, -- in t_slv_8_arr(1 downto 0);
--        data2_i => data2, -- in t_slv_8_arr(1 downto 0);
--        data3_i => data3, -- in t_slv_8_arr(1 downto 0);
--        meta_i  => correlatorMetaIn, -- in std_logic_vector((METABITS-1) downto 0);  -- Sampled on the first cycle of every third packet of valid_i. 
--        valid_i => DataValid,    -- in std_logic;
--        -- Data out; bursts of 216 clocks for each channel.
--        data0_o => corFBDout0,    -- out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
--        data1_o => corFBDout1,    -- out t_slv_16_arr(1 downto 0);
--        data2_o => corFBDout2,    -- out t_slv_16_arr(1 downto 0);
--        data3_o => corFBDout3,    -- out t_slv_16_arr(1 downto 0);
        
--        meta_o  => corMetaOut,  -- out std_logic_vector((METABITS-1) downto 0);
--        valid_o => corValidOut, -- out std_logic;
--        -- Writing FIR Taps
--        FIRTapData_i   => (others => '0'),  -- in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
--        FIRTapData_o   => open,             -- out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
--        FIRTapAddr_i   => (others => '0'),  -- in std_logic_vector(15 downto 0);   -- 4096 * 12 filter taps = 49152 total.
--        FIRTapWE_i     => '0',              -- in std_logic;
--        FIRTapClk      => i_axi_clk         -- in std_logic;
--    );
    
    corfbi : entity filterbanks_lib.correlatorFBTop_dummy
    generic map(
        METABITS => 620,    -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP => 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    ) port map (
        -- clock, target is 380 MHz
        clk  => i_axi_clk, -- in std_logic;
        rst  => i_SOF,     -- in std_logic;
        -- Data input, common valid signal, expects packets of 4096 samples. Requires at least 2 clocks idle time between packets.
        meta_i  => correlatorMetaIn,
        valid_i => DataValid,
        
        -- Data out; bursts of 3456 clocks for each channel.
        meta_o  => corMetaOut,  -- out std_logic_vector((METABITS-1) downto 0);
        valid_o => corValidOut
    );
    
    
--    corfb2i : entity filterbanks_lib.correlatorFBTop25
--    generic map(
--        METABITS => 361,    -- Width in bits of the meta_i and meta_o ports.
--        FRAMESTODROP => 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
--    ) port map (
--        -- processing clock
--        clk     => i_axi_clk,
--        rst     => i_SOF,
--        -- Data input, common valid signal, expects packets of 64 samples. 
--        -- Requires at least 2 clocks idle time between packets.
--        -- Due to oversampling, also requires on average 86 clocks between packets - specifically, no more than 3 packets in 258 clocks. 
--        data0_i => data4, -- in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
--        data1_i => data5, -- in t_slv_8_arr(1 downto 0);
--        data2_i => data6, -- in t_slv_8_arr(1 downto 0);
--        data3_i => data7, -- in t_slv_8_arr(1 downto 0);
--        meta_i  => correlatorMetaIn, -- in std_logic_vector((METABITS-1) downto 0);  -- Sampled on the first cycle of every third packet of valid_i. 
--        valid_i => DataValid,    -- in std_logic;
--        -- Data out; bursts of 216 clocks for each channel.
--        data0_o => corFBDout4,    -- out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
--        data1_o => corFBDout5,    -- out t_slv_16_arr(1 downto 0);
--        data2_o => corFBDout6,    -- out t_slv_16_arr(1 downto 0);
--        data3_o => corFBDout7,    -- out t_slv_16_arr(1 downto 0);
        
--        meta_o  => open,  -- out std_logic_vector((METABITS-1) downto 0);
--        valid_o => open,  -- out std_logic;
--        -- Writing FIR Taps
--        FIRTapData_i   => (others => '0'),  -- in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
--        FIRTapData_o   => open,             -- out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
--        FIRTapAddr_i   => (others => '0'),  -- in std_logic_vector(15 downto 0);   -- 4096 * 12 filter taps = 49152 total.
--        FIRTapWE_i     => '0',              -- in std_logic;
--        FIRTapClk      => i_axi_clk         -- in std_logic;
--    );
    
    -- Pack the filterbank output into a structure for input to the fine delay module.
    corDout_arr(0).vpol.re <= corFBDout0(0);  -- 16 bit data into the fine delay module.
    corDout_arr(0).vpol.im <= corFBDout0(1);
    corDout_arr(0).hpol.re <= corFBDout1(0);
    corDout_arr(0).hpol.im <= corFBDout1(1);
    corDout_arr(1).vpol.re <= corFBDout2(0);  -- 16 bit data into the fine delay module.
    corDout_arr(1).vpol.im <= corFBDout2(1);
    corDout_arr(1).hpol.re <= corFBDout3(0);
    corDout_arr(1).hpol.im <= corFBDout3(1);
    corDout_arr(2).vpol.re <= corFBDout4(0);  -- 16 bit data into the fine delay module.
    corDout_arr(2).vpol.im <= corFBDout4(1);
    corDout_arr(2).hpol.re <= corFBDout5(0);
    corDout_arr(2).hpol.im <= corFBDout5(1);
    corDout_arr(3).vpol.re <= corFBDout6(0);  -- 16 bit data into the fine delay module.
    corDout_arr(3).vpol.im <= corFBDout6(1);
    corDout_arr(3).hpol.re <= corFBDout7(0);
    corDout_arr(3).hpol.im <= corFBDout7(1);
    
    --o_CorDataValid <= CorValidOut;
    corFBHeader(0).HDeltaP          <= corMetaOut(31 downto 0);
    corFBHeader(0).VDeltaP          <= corMetaOut(63 downto 32);
    corFBHeader(0).HOffsetP         <= corMetaOut(95 downto 64);
    corFBHeader(0).VOffsetP         <= corMetaOut(127 downto 96);
    corFBHeader(0).virtualChannel   <= corMetaOut(143 downto 128);
    corFBHeader(0).valid            <= corMetaOut(144);
    corFBHeader(0).integration      <= corMetaOut(31+580 downto 0+580);
    corFBHeader(0).ctFrame          <= corMetaOut(33+580 downto 32+580);
    corFBHeader(0).bad_poly <= corMetaOut(614);
    corFBHeader(0).lastChannel <= corMetaOut(618);
    corFBHeader(0).demap_table_select <= corMetaOut(619);
    
    corFBHeader(1).HDeltaP          <= corMetaOut(31+145 downto 0+145);
    corFBHeader(1).VDeltaP          <= corMetaOut(63+145 downto 32+145);
    corFBHeader(1).HOffsetP         <= corMetaOut(95+145 downto 64+145);
    corFBHeader(1).VOffsetP         <= corMetaOut(127+145 downto 96+145);
    corFBHeader(1).virtualChannel   <= corMetaOut(143+145 downto 128+145);
    corFBHeader(1).valid            <= corMetaOut(144+145);
    corFBHeader(1).integration      <= corMetaOut(31+580 downto 0+580);
    corFBHeader(1).ctFrame          <= corMetaOut(33+580 downto 32+580);
    corFBHeader(1).bad_poly <= corMetaOut(615);
    corFBHeader(1).lastChannel <= corMetaOut(618);
    corFBHeader(1).demap_table_select <= corMetaOut(619);
    
    corFBHeader(2).HDeltaP          <= corMetaOut(31+290 downto 0+290);
    corFBHeader(2).VDeltaP          <= corMetaOut(63+290 downto 32+290);
    corFBHeader(2).HOffsetP         <= corMetaOut(95+290 downto 64+290);
    corFBHeader(2).VOffsetP         <= corMetaOut(127+290 downto 96+290);
    corFBHeader(2).virtualChannel   <= corMetaOut(143+290 downto 128+290);
    corFBHeader(2).valid            <= corMetaOut(144+290);
    corFBHeader(2).integration      <= corMetaOut(31+580 downto 0+580);
    corFBHeader(2).ctFrame          <= corMetaOut(33+580 downto 32+580);
    corFBHeader(2).bad_poly <= corMetaOut(616);
    corFBHeader(2).lastChannel <= corMetaOut(618);
    corFBHeader(2).demap_table_select <= corMetaOut(619);
    
    corFBHeader(3).HDeltaP          <= corMetaOut(31+435 downto 0+435);
    corFBHeader(3).VDeltaP          <= corMetaOut(63+435 downto 32+435);
    corFBHeader(3).HOffsetP         <= corMetaOut(95+435 downto 64+435);
    corFBHeader(3).VOffsetP         <= corMetaOut(127+435 downto 96+435);
    corFBHeader(3).virtualChannel   <= corMetaOut(143+435 downto 128+435);
    corFBHeader(3).valid            <= corMetaOut(144+435);
    corFBHeader(3).integration      <= corMetaOut(31+580 downto 0+580);
    corFBHeader(3).ctFrame          <= corMetaOut(33+580 downto 32+580);
    corFBHeader(3).bad_poly <= corMetaOut(617);
    corFBHeader(3).lastChannel <= corMetaOut(618);
    corFBHeader(3).demap_table_select <= corMetaOut(619);
    
    corFBHeaderValid <= corValidOut and (not corValidOutDel);
    
    process(i_axi_clk)
    begin
        if rising_edge(i_axi_clk) then
            corValidOutDel <= corValidOut;
        end if;
    end process;
    
--    FDGen : for i in 0 to 3 generate 
--        FineDelay : entity filterbanks_lib.fineDelay
--        generic map (
--            FBSELECTION => 2  -- 2 = Correlator
--        )
--        port map (
--            i_clk  => i_axi_clk,
--            -- data and header in
--            i_data        => corDout_arr(i),    --  in t_FB_output_payload;  -- 16 bit data : .Hpol.re, Hpol.im, .Vpol.re, .Vpol.im 
--            i_dataValid   => corValidOut,       -- in std_logic;
--            i_header      => corFBHeader(i),    -- in t_atomic_CT_pst_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(36:0), virtualChannel(15:0), .valid
--            i_headerValid => corFBHeaderValid,  -- in std_logic;
--            -- Data and Header out
--            o_data        => FDdata(i),         -- out t_ctc_output_payload;   -- 8 bit data : .Hpol.re, Hpol.im, .Vpol.re, .Vpol.im 
--            o_dataValid   => FDcorDataValid(i), -- out std_logic;
--            o_header      => FDHeader(i),       -- out t_atomic_CT_pst_META_out; -- .HDeltaP(15:0), .VDeltaP(15:0), .frameCount(36:0), virtualChannel(15:0), .valid
--            o_headerValid => headerValid(i),    -- out std_logic;
    
--            -------------------------------------------
--            -- control and monitoring
--            -- Disable the fine delay. Instead of multiplying by the output of the sin/cos lookup, just scale by unity.
--            i_disable     => i_fineDelayDisable, -- in std_logic;
--            -- Scale down by 2^(i_RFIScale) before clipping for RFI.
--            -- Unity for the sin/cos lookup is 0x10000, so :
--            --   i_RFIScale < 16  ==> Amplify the output of the filterbanks.
--            --   i_RFIScale = 16  ==> Amplitude of the filterbank output is unchanged.
--            --   i_RFIScale > 16  ==> Amplitude of the filterbank output is reduced.
--            i_RFIScale    => i_RFIScale, -- in std_logic_vector(4 downto 0); 
--            -- For monitoring of the output level.
--            -- Higher level should keep track of : 
--            --   * The total number of frames processed.
--            --   * The sum of each of the outputs below. (but note one is superfluous since it can be calculated from the total frames processed and the sum of all the others).
--            --      - These sums should be 32 bit values, which ensures wrapping will occur at most once per hour.
--            -- For the correlator:
--            --   - Each frame corresponds to 3456 fine channels x 2 (H & V polarisations) * 2 (re+im).
--            --   - Every fine channel must be one of the categories below, so they will sum to 3456*2*2 = 13824.
--            o_overflow    => open, -- hist_overflow(i),     -- out(15:0); -- Number of fine channels which were clipped.
--            o_64_127      => open, -- hist_64_127(i),  -- out(15:0); -- Number of fine channels in the range 64 to 128.
--            o_32_63       => open, -- hist_32_63(i),   -- out(15:0); -- Number of fine channels in the range 32 to 64.
--            o_16_31       => open, -- hist_16_31(i),   -- out(15:0); -- Number of fine channels in the range 16 to 32.
--            o_0_15        => open, -- hist_0_15(i),    -- out(15:0); -- Number of fine channels in the range 0 to 15.
--            o_virtualChannel => open, -- hist_virtualChannel(i), -- out(8:0);
--            o_histogramValid => open  -- hist_valid(i) -- out std_logic -- indicates histogram data is valid.
--        );
--    end generate;
    
    -- fineDelay incurs a 19 clock latency on the data.
    process(i_axi_clk)
    begin
        if rising_edge(i_axi_clk) then
            FD_virtualChannel0(0) <= corFBHeader(0).virtualChannel(15 downto 0);
            FD_virtualChannel0(18 downto 1) <= FD_virtualChannel0(17 downto 0);
            FD_virtualChannel1(0) <= corFBHeader(1).virtualChannel(15 downto 0);
            FD_virtualChannel1(18 downto 1) <= FD_virtualChannel1(17 downto 0);
            FD_virtualChannel2(0) <= corFBHeader(2).virtualChannel(15 downto 0);
            FD_virtualChannel2(18 downto 1) <= FD_virtualChannel2(17 downto 0);
            FD_virtualChannel3(0) <= corFBHeader(3).virtualChannel(15 downto 0);
            FD_virtualChannel3(18 downto 1) <= FD_virtualChannel3(17 downto 0);
            
            FD_bad_poly(0) <= corFBHeader(0).bad_poly or corFBHeader(1).bad_poly or corFBHeader(2).bad_poly or corFBHeader(3).bad_poly;
            FD_bad_poly(18 downto 1) <= FD_bad_poly(17 downto 0);
            
            FD_lastChannel(0) <= corFBHeader(0).lastChannel;
            FD_lastChannel(18 downto 1) <= FD_lastChannel(17 downto 0);
            FD_demap_table_select(0) <= corFBHeader(0).demap_table_select;
            FD_demap_table_select(18 downto 1) <= FD_demap_table_select(17 downto 0);
            
            FD_integration(0) <= corFBHeader(0).integration;
            FD_integration(18 downto 1) <= FD_integration(17 downto 0);
            
            FD_ctFrame(0) <= corFBHeader(0).ctFrame;
            FD_ctFrame(18 downto 1) <= FD_ctFrame(17 downto 0);
             
            FD_datavalid(0) <= corValidOut;
            FD_datavalid(18 downto 1) <= FD_datavalid(17 downto 0);
            
            FD_headerValid(0) <= corFBHeaderValid;
            FD_headerValid(18 downto 1) <= FD_headerValid(17 downto 0);
            
            if FD_datavalid(18) = '0' then
                FD_finecount <= x"0000";
            else
                FD_finecount <= std_logic_vector(unsigned(FD_finecount) + 1);
            end if;
        end if;
    end process;
        
    o_data(0).Hpol.re <= FD_virtualChannel0(18)(7 downto 0);
    o_data(0).Hpol.im <= FD_integration(18)(7 downto 0);
    o_data(0).Vpol.re <= FD_finecount(7 downto 0);
    o_data(0).Vpol.im <= FD_finecount(15 downto 8);

    o_data(1).Hpol.re <= FD_virtualChannel1(18)(7 downto 0);
    o_data(1).Hpol.im <= FD_integration(18)(7 downto 0);
    o_data(1).Vpol.re <= FD_finecount(7 downto 0);
    o_data(1).Vpol.im <= FD_finecount(15 downto 8);
    
    o_data(2).Hpol.re <= FD_virtualChannel2(18)(7 downto 0);
    o_data(2).Hpol.im <= FD_integration(18)(7 downto 0);
    o_data(2).Vpol.re <= FD_finecount(7 downto 0);
    o_data(2).Vpol.im <= FD_finecount(15 downto 8);
    
    o_data(3).Hpol.re <= FD_virtualChannel3(18)(7 downto 0);
    o_data(3).Hpol.im <= FD_integration(18)(7 downto 0);
    o_data(3).Vpol.re <= FD_finecount(7 downto 0);
    o_data(3).Vpol.im <= FD_finecount(15 downto 8);
    
    o_dataValid <= FD_datavalid(18);
    o_virtualChannel(0) <= FD_virtualChannel0(18);
    o_virtualChannel(1) <= FD_virtualChannel1(18);
    o_virtualChannel(2) <= FD_virtualChannel2(18);
    o_virtualChannel(3) <= FD_virtualChannel3(18);
    o_bad_poly <= FD_bad_poly(18);
    o_lastChannel <= FD_lastChannel(18);
    o_demap_table_select <= FD_demap_table_select(18);
    
    o_integration <= FD_integration(18);
    o_ctFrame <= FD_ctFrame(18);
    o_headerValid(0) <= FD_headerValid(18);
    o_headerValid(1) <= FD_headerValid(18);
    o_headerValid(2) <= FD_headerValid(18);
    o_headerValid(3) <= FD_headerValid(18);
    
--    o_data <= FDdata;
--    o_dataValid <= FDcorDataValid(0);  -- FDPSTDataValid(0) and (1), (2), (3) will be the same.
--    o_virtualChannel(0) <= FDHeader(0).virtualChannel;
--    o_virtualChannel(1) <= FDHeader(1).virtualChannel;
--    o_virtualChannel(2) <= FDHeader(2).virtualChannel;
--    o_virtualChannel(3) <= FDHeader(3).virtualChannel;
--    o_frameCount <= FDHeader(0).frameCount;
--    o_headerValid <= headerValid;
    ---------------------------------------------------------------
    -- Registers
    -- 
    
    filterbank_Reg : entity filterbanks_lib.cor_filterbanks_filterbanks_reg
    port map(
        MM_CLK              => i_axi_clk,   -- in  std_logic;
        MM_RST              => i_axi_rst,   -- in  std_logic;
        SLA_IN              => i_axi_mosi,  -- IN  t_axi4_lite_mosi;
        SLA_OUT             => o_axi_miso,  -- OUT t_axi4_lite_miso;
        CONFIG_FIELDS_RO	=> config_ro,   -- IN  t_config_ro;
        CONFIG_FIELDS_RW    => config_rw,   -- out t_config_rw;
        CONFIG_OUTPUT_DISABLE_IN  => output_disable_i, -- IN  t_config_output_disable_ram_in;
        CONFIG_OUTPUT_DISABLE_OUT => output_disable_o  -- OUT t_config_output_disable_ram_out
    );
    
    config_ro.status <= x"00000000";
    config_ro.txCount_eth <= tx_packet_count;
    config_ro.txcount_corner_turn <= tx_packet_count_ct;
    
    process(i_axi_clk)
    begin
        if rising_edge(i_axi_clk) then
            reg_reset <= config_rw.config(0);
            reg_reset_del1 <= reg_reset;
            
            -- count of ethernet packet going out.
            if reg_reset = '1' and reg_reset_del1 = '0' then
                tx_packet_count <= (others => '0');
            elsif packetValid = '1' and packetValidDel1 = '0' then
                tx_packet_count <= std_logic_vector(unsigned(tx_packet_count) + 1);
            end if;
            
            -- count of packets going out to the corner turn.
            FDcorDataValidDel <= FDcorDataValid(0);
            if reg_reset = '1' and reg_reset_del1 = '0' then
                tx_packet_count_ct <= (others => '0');
            elsif FDcorDataValid(0) = '1' and FDcorDataValidDel = '0' then
                tx_packet_count_ct <= std_logic_vector(unsigned(tx_packet_count_ct) + 1);
            end if;
            
        end if;
    end process;
    
    output_disable_i.adr <= output_disable_addr;
    output_disable_i.wr_dat <= (others => '0');
    output_disable_i.wr_en <= '0';
    output_disable_i.rd_en <= '1';
    output_disable_i.clk <= i_axi_clk;
    output_disable_i.rst <= '0';
    
    --------------------------------------------------------------
    -- Packets of samples to go to the 100G
    -- Each output packet contains : 
    --  16 byte header : 
    --    5 bytes = 40 bits : framecount
    --    2 bytes = 16 bits : virtual channel
    --    1 byte  = 8  bits : Polarisation (either 0 or 1)
    --    8 bytes           : unused.
    --  Data : 
    --    8+8 bit complex data for 3456 fine channels.
    --    = 6912 bytes of data.
    
    -- Buffer : The output from the fine delay arrives as a burst, with
    --  16 bytes wide; 3456 clocks long.
    -- This double buffers the data so that we can output packets with data for a single
    -- coarse channel and polarisation in a single packet.
    -- The buffer is split into 16 x (512 deep) pages, 2 buffers for each of
    --  coarse 0, pol 0, 
    --  coarse 0, pol 1,
    --  coarse 1, pol 0,
    --  coarse 1, pol 1,
    --  coarse 2, pol 0, 
    --  coarse 2, pol 1,
    --  coarse 3, pol 0, 
    --  coarse 3, pol 1,
    
    o_packetValid <= '0';
    o_packetData <= (others => '0');
    
    
    
end Behavioral;