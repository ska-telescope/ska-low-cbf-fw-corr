-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom5 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom5; 
 
architecture behavioral of inv_rom5 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"39cccccd", 
    x"39ccb854", 
    x"39cca3df", 
    x"39cc8f6f", 
    x"39cc7b02", 
    x"39cc669a", 
    x"39cc5235", 
    x"39cc3dd5", 
    x"39cc2978", 
    x"39cc1520", 
    x"39cc00cc", 
    x"39cbec7c", 
    x"39cbd830", 
    x"39cbc3e8", 
    x"39cbafa4", 
    x"39cb9b64", 
    x"39cb8728", 
    x"39cb72f0", 
    x"39cb5ebc", 
    x"39cb4a8c", 
    x"39cb3660", 
    x"39cb2238", 
    x"39cb0e14", 
    x"39caf9f4", 
    x"39cae5d8", 
    x"39cad1c0", 
    x"39cabdac", 
    x"39caa99c", 
    x"39ca9590", 
    x"39ca8188", 
    x"39ca6d84", 
    x"39ca5984", 
    x"39ca4588", 
    x"39ca3190", 
    x"39ca1d9b", 
    x"39ca09ab", 
    x"39c9f5bf", 
    x"39c9e1d6", 
    x"39c9cdf1", 
    x"39c9ba11", 
    x"39c9a634", 
    x"39c9925b", 
    x"39c97e86", 
    x"39c96ab5", 
    x"39c956e8", 
    x"39c9431f", 
    x"39c92f59", 
    x"39c91b98", 
    x"39c907da", 
    x"39c8f421", 
    x"39c8e06b", 
    x"39c8ccb9", 
    x"39c8b90b", 
    x"39c8a560", 
    x"39c891ba", 
    x"39c87e17", 
    x"39c86a79", 
    x"39c856de", 
    x"39c84347", 
    x"39c82fb3", 
    x"39c81c24", 
    x"39c80898", 
    x"39c7f511", 
    x"39c7e18d", 
    x"39c7ce0c", 
    x"39c7ba90", 
    x"39c7a718", 
    x"39c793a3", 
    x"39c78032", 
    x"39c76cc5", 
    x"39c7595b", 
    x"39c745f6", 
    x"39c73294", 
    x"39c71f36", 
    x"39c70bdb", 
    x"39c6f885", 
    x"39c6e532", 
    x"39c6d1e3", 
    x"39c6be98", 
    x"39c6ab50", 
    x"39c6980c", 
    x"39c684cc", 
    x"39c67190", 
    x"39c65e57", 
    x"39c64b22", 
    x"39c637f1", 
    x"39c624c4", 
    x"39c6119a", 
    x"39c5fe74", 
    x"39c5eb52", 
    x"39c5d833", 
    x"39c5c518", 
    x"39c5b201", 
    x"39c59eed", 
    x"39c58bdd", 
    x"39c578d1", 
    x"39c565c8", 
    x"39c552c4", 
    x"39c53fc2", 
    x"39c52cc5", 
    x"39c519cb", 
    x"39c506d5", 
    x"39c4f3e2", 
    x"39c4e0f3", 
    x"39c4ce08", 
    x"39c4bb20", 
    x"39c4a83c", 
    x"39c4955b", 
    x"39c4827f", 
    x"39c46fa5", 
    x"39c45cd0", 
    x"39c449fe", 
    x"39c43730", 
    x"39c42465", 
    x"39c4119e", 
    x"39c3feda", 
    x"39c3ec1a", 
    x"39c3d95e", 
    x"39c3c6a5", 
    x"39c3b3f0", 
    x"39c3a13e", 
    x"39c38e90", 
    x"39c37be5", 
    x"39c3693e", 
    x"39c3569b", 
    x"39c343fb", 
    x"39c3315f", 
    x"39c31ec6", 
    x"39c30c31", 
    x"39c2f99f", 
    x"39c2e711", 
    x"39c2d486", 
    x"39c2c1ff", 
    x"39c2af7c", 
    x"39c29cfc", 
    x"39c28a7f", 
    x"39c27806", 
    x"39c26591", 
    x"39c2531f", 
    x"39c240b0", 
    x"39c22e45", 
    x"39c21bde", 
    x"39c20979", 
    x"39c1f719", 
    x"39c1e4bc", 
    x"39c1d262", 
    x"39c1c00c", 
    x"39c1adb9", 
    x"39c19b6a", 
    x"39c1891f", 
    x"39c176d6", 
    x"39c16491", 
    x"39c15250", 
    x"39c14012", 
    x"39c12dd8", 
    x"39c11ba1", 
    x"39c1096d", 
    x"39c0f73d", 
    x"39c0e510", 
    x"39c0d2e7", 
    x"39c0c0c1", 
    x"39c0ae9e", 
    x"39c09c7f", 
    x"39c08a63", 
    x"39c0784b", 
    x"39c06636", 
    x"39c05425", 
    x"39c04217", 
    x"39c0300c", 
    x"39c01e05", 
    x"39c00c01", 
    x"39bffa00", 
    x"39bfe803", 
    x"39bfd609", 
    x"39bfc413", 
    x"39bfb220", 
    x"39bfa030", 
    x"39bf8e44", 
    x"39bf7c5b", 
    x"39bf6a75", 
    x"39bf5892", 
    x"39bf46b4", 
    x"39bf34d8", 
    x"39bf2300", 
    x"39bf112b", 
    x"39beff59", 
    x"39beed8b", 
    x"39bedbc0", 
    x"39bec9f8", 
    x"39beb833", 
    x"39bea672", 
    x"39be94b5", 
    x"39be82fa", 
    x"39be7143", 
    x"39be5f8f", 
    x"39be4dde", 
    x"39be3c31", 
    x"39be2a87", 
    x"39be18e0", 
    x"39be073d", 
    x"39bdf59d", 
    x"39bde400", 
    x"39bdd266", 
    x"39bdc0d0", 
    x"39bdaf3c", 
    x"39bd9dac", 
    x"39bd8c20", 
    x"39bd7a96", 
    x"39bd6910", 
    x"39bd578d", 
    x"39bd460e", 
    x"39bd3491", 
    x"39bd2318", 
    x"39bd11a2", 
    x"39bd002f", 
    x"39bceec0", 
    x"39bcdd53", 
    x"39bccbea", 
    x"39bcba84", 
    x"39bca922", 
    x"39bc97c2", 
    x"39bc8666", 
    x"39bc750d", 
    x"39bc63b7", 
    x"39bc5264", 
    x"39bc4114", 
    x"39bc2fc8", 
    x"39bc1e7f", 
    x"39bc0d39", 
    x"39bbfbf6", 
    x"39bbeab6", 
    x"39bbd97a", 
    x"39bbc841", 
    x"39bbb70a", 
    x"39bba5d7", 
    x"39bb94a7", 
    x"39bb837b", 
    x"39bb7251", 
    x"39bb612b", 
    x"39bb5007", 
    x"39bb3ee7", 
    x"39bb2dca", 
    x"39bb1cb0", 
    x"39bb0b99", 
    x"39bafa86", 
    x"39bae975", 
    x"39bad868", 
    x"39bac75d", 
    x"39bab656", 
    x"39baa552", 
    x"39ba9451", 
    x"39ba8353", 
    x"39ba7258", 
    x"39ba6160", 
    x"39ba506c", 
    x"39ba3f7a", 
    x"39ba2e8c", 
    x"39ba1da0", 
    x"39ba0cb8", 
    x"39b9fbd3", 
    x"39b9eaf0", 
    x"39b9da11", 
    x"39b9c935", 
    x"39b9b85c", 
    x"39b9a786", 
    x"39b996b3", 
    x"39b985e3", 
    x"39b97517", 
    x"39b9644d", 
    x"39b95386", 
    x"39b942c2", 
    x"39b93202", 
    x"39b92144", 
    x"39b91089", 
    x"39b8ffd2", 
    x"39b8ef1d", 
    x"39b8de6c", 
    x"39b8cdbd", 
    x"39b8bd11", 
    x"39b8ac69", 
    x"39b89bc3", 
    x"39b88b21", 
    x"39b87a81", 
    x"39b869e5", 
    x"39b8594b", 
    x"39b848b5", 
    x"39b83821", 
    x"39b82791", 
    x"39b81703", 
    x"39b80678", 
    x"39b7f5f1", 
    x"39b7e56c", 
    x"39b7d4ea", 
    x"39b7c46b", 
    x"39b7b3ef", 
    x"39b7a377", 
    x"39b79301", 
    x"39b7828e", 
    x"39b7721e", 
    x"39b761b1", 
    x"39b75147", 
    x"39b740df", 
    x"39b7307b", 
    x"39b7201a", 
    x"39b70fbb", 
    x"39b6ff60", 
    x"39b6ef07", 
    x"39b6deb2", 
    x"39b6ce5f", 
    x"39b6be0f", 
    x"39b6adc2", 
    x"39b69d78", 
    x"39b68d31", 
    x"39b67ced", 
    x"39b66cac", 
    x"39b65c6d", 
    x"39b64c32", 
    x"39b63bf9", 
    x"39b62bc4", 
    x"39b61b91", 
    x"39b60b61", 
    x"39b5fb34", 
    x"39b5eb09", 
    x"39b5dae2", 
    x"39b5cabe", 
    x"39b5ba9c", 
    x"39b5aa7d", 
    x"39b59a61", 
    x"39b58a48", 
    x"39b57a32", 
    x"39b56a1f", 
    x"39b55a0e", 
    x"39b54a01", 
    x"39b539f6", 
    x"39b529ee", 
    x"39b519e9", 
    x"39b509e7", 
    x"39b4f9e7", 
    x"39b4e9ea", 
    x"39b4d9f1", 
    x"39b4c9fa", 
    x"39b4ba05", 
    x"39b4aa14", 
    x"39b49a26", 
    x"39b48a3a", 
    x"39b47a51", 
    x"39b46a6b", 
    x"39b45a87", 
    x"39b44aa7", 
    x"39b43ac9", 
    x"39b42aee", 
    x"39b41b16", 
    x"39b40b41", 
    x"39b3fb6e", 
    x"39b3eb9e", 
    x"39b3dbd1", 
    x"39b3cc07", 
    x"39b3bc40", 
    x"39b3ac7b", 
    x"39b39cb9", 
    x"39b38cfa", 
    x"39b37d3d", 
    x"39b36d84", 
    x"39b35dcd", 
    x"39b34e19", 
    x"39b33e67", 
    x"39b32eb8", 
    x"39b31f0d", 
    x"39b30f63", 
    x"39b2ffbd", 
    x"39b2f019", 
    x"39b2e078", 
    x"39b2d0da", 
    x"39b2c13e", 
    x"39b2b1a6", 
    x"39b2a210", 
    x"39b2927c", 
    x"39b282ec", 
    x"39b2735e", 
    x"39b263d2", 
    x"39b2544a", 
    x"39b244c4", 
    x"39b23541", 
    x"39b225c1", 
    x"39b21643", 
    x"39b206c8", 
    x"39b1f74f", 
    x"39b1e7da", 
    x"39b1d867", 
    x"39b1c8f7", 
    x"39b1b989", 
    x"39b1aa1e", 
    x"39b19ab6", 
    x"39b18b50", 
    x"39b17bed", 
    x"39b16c8d", 
    x"39b15d2f", 
    x"39b14dd5", 
    x"39b13e7c", 
    x"39b12f27", 
    x"39b11fd4", 
    x"39b11083", 
    x"39b10136", 
    x"39b0f1eb", 
    x"39b0e2a2", 
    x"39b0d35d", 
    x"39b0c41a", 
    x"39b0b4d9", 
    x"39b0a59b", 
    x"39b09660", 
    x"39b08727", 
    x"39b077f2", 
    x"39b068be", 
    x"39b0598d", 
    x"39b04a5f", 
    x"39b03b34", 
    x"39b02c0b", 
    x"39b01ce5", 
    x"39b00dc1", 
    x"39affea0", 
    x"39afef82", 
    x"39afe066", 
    x"39afd14c", 
    x"39afc236", 
    x"39afb322", 
    x"39afa410", 
    x"39af9501", 
    x"39af85f5", 
    x"39af76eb", 
    x"39af67e4", 
    x"39af58df", 
    x"39af49dd", 
    x"39af3ade", 
    x"39af2be1", 
    x"39af1ce7", 
    x"39af0def", 
    x"39aefefa", 
    x"39aef007", 
    x"39aee117", 
    x"39aed229", 
    x"39aec33e", 
    x"39aeb456", 
    x"39aea570", 
    x"39ae968c", 
    x"39ae87ab", 
    x"39ae78cd", 
    x"39ae69f1", 
    x"39ae5b18", 
    x"39ae4c41", 
    x"39ae3d6d", 
    x"39ae2e9b", 
    x"39ae1fcc", 
    x"39ae1100", 
    x"39ae0236", 
    x"39adf36e", 
    x"39ade4a9", 
    x"39add5e6", 
    x"39adc726", 
    x"39adb869", 
    x"39ada9ad", 
    x"39ad9af5", 
    x"39ad8c3f", 
    x"39ad7d8b", 
    x"39ad6eda", 
    x"39ad602b", 
    x"39ad517f", 
    x"39ad42d6", 
    x"39ad342e", 
    x"39ad258a", 
    x"39ad16e7", 
    x"39ad0848", 
    x"39acf9aa", 
    x"39aceb10", 
    x"39acdc77", 
    x"39accde1", 
    x"39acbf4e", 
    x"39acb0bd", 
    x"39aca22e", 
    x"39ac93a2", 
    x"39ac8519", 
    x"39ac7692", 
    x"39ac680d", 
    x"39ac598b", 
    x"39ac4b0b", 
    x"39ac3c8d", 
    x"39ac2e12", 
    x"39ac1f9a", 
    x"39ac1124", 
    x"39ac02b0", 
    x"39abf43f", 
    x"39abe5d0", 
    x"39abd764", 
    x"39abc8fa", 
    x"39abba92", 
    x"39abac2d", 
    x"39ab9dca", 
    x"39ab8f6a", 
    x"39ab810c", 
    x"39ab72b0", 
    x"39ab6457", 
    x"39ab5601", 
    x"39ab47ac", 
    x"39ab395a", 
    x"39ab2b0b", 
    x"39ab1cbe", 
    x"39ab0e73", 
    x"39ab002b", 
    x"39aaf1e5", 
    x"39aae3a1", 
    x"39aad560", 
    x"39aac721", 
    x"39aab8e5"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
