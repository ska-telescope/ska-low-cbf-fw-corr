-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom0 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom0; 
 
architecture behavioral of inv_rom0 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"3b004020", 
    x"3b008081", 
    x"3b00c122", 
    x"3b010204", 
    x"3b014328", 
    x"3b01848e", 
    x"3b01c636", 
    x"3b020821", 
    x"3b024a4e", 
    x"3b028cc0", 
    x"3b02cf75", 
    x"3b03126f", 
    x"3b0355ad", 
    x"3b039930", 
    x"3b03dcf9", 
    x"3b042108", 
    x"3b04655e", 
    x"3b04a9fa", 
    x"3b04eedd", 
    x"3b053408", 
    x"3b05797c", 
    x"3b05bf37", 
    x"3b06053c", 
    x"3b064b8a", 
    x"3b069223", 
    x"3b06d905", 
    x"3b072033", 
    x"3b0767ab", 
    x"3b07af70", 
    x"3b07f781", 
    x"3b083fde", 
    x"3b088889", 
    x"3b08d181", 
    x"3b091ac7", 
    x"3b09645c", 
    x"3b09ae41", 
    x"3b09f874", 
    x"3b0a42f8", 
    x"3b0a8dcd", 
    x"3b0ad8f3", 
    x"3b0b246b", 
    x"3b0b7034", 
    x"3b0bbc51", 
    x"3b0c08c1", 
    x"3b0c5584", 
    x"3b0ca29c", 
    x"3b0cf009", 
    x"3b0d3dcb", 
    x"3b0d8be3", 
    x"3b0dda52", 
    x"3b0e2918", 
    x"3b0e7835", 
    x"3b0ec7ab", 
    x"3b0f177a", 
    x"3b0f67a2", 
    x"3b0fb824", 
    x"3b100901", 
    x"3b105a38", 
    x"3b10abcc", 
    x"3b10fdbc", 
    x"3b115009", 
    x"3b11a2b4", 
    x"3b11f5bd", 
    x"3b124925", 
    x"3b129cec", 
    x"3b12f114", 
    x"3b13459c", 
    x"3b139a86", 
    x"3b13efd2", 
    x"3b144581", 
    x"3b149b93", 
    x"3b14f209", 
    x"3b1548e5", 
    x"3b15a025", 
    x"3b15f7cc", 
    x"3b164fda", 
    x"3b16a850", 
    x"3b17012e", 
    x"3b175a75", 
    x"3b17b426", 
    x"3b180e41", 
    x"3b1868c8", 
    x"3b18c3bb", 
    x"3b191f1a", 
    x"3b197ae7", 
    x"3b19d723", 
    x"3b1a33cd", 
    x"3b1a90e8", 
    x"3b1aee73", 
    x"3b1b4c70", 
    x"3b1baadf", 
    x"3b1c09c1", 
    x"3b1c6917", 
    x"3b1cc8e1", 
    x"3b1d2922", 
    x"3b1d89d9", 
    x"3b1deb07", 
    x"3b1e4cad", 
    x"3b1eaecd", 
    x"3b1f1166", 
    x"3b1f747a", 
    x"3b1fd80a", 
    x"3b203c17", 
    x"3b20a0a1", 
    x"3b2105a9", 
    x"3b216b31", 
    x"3b21d13a", 
    x"3b2237c3", 
    x"3b229ecf", 
    x"3b23065e", 
    x"3b236e72", 
    x"3b23d70a", 
    x"3b244029", 
    x"3b24a9cf", 
    x"3b2513fd", 
    x"3b257eb5", 
    x"3b25e9f7", 
    x"3b2655c4", 
    x"3b26c21e", 
    x"3b272f05", 
    x"3b279c7b", 
    x"3b280a81", 
    x"3b287917", 
    x"3b28e83f", 
    x"3b2957fb", 
    x"3b29c84a", 
    x"3b2a392f", 
    x"3b2aaaab", 
    x"3b2b1cbe", 
    x"3b2b8f6a", 
    x"3b2c02b0", 
    x"3b2c7692", 
    x"3b2ceb10", 
    x"3b2d602b", 
    x"3b2dd5e6", 
    x"3b2e4c41", 
    x"3b2ec33e", 
    x"3b2f3ade", 
    x"3b2fb322", 
    x"3b302c0b", 
    x"3b30a59b", 
    x"3b311fd4", 
    x"3b319ab6", 
    x"3b321643", 
    x"3b32927c", 
    x"3b330f63", 
    x"3b338cfa", 
    x"3b340b41", 
    x"3b348a3a", 
    x"3b3509e7", 
    x"3b358a48", 
    x"3b360b61", 
    x"3b368d31", 
    x"3b370fbb", 
    x"3b379301", 
    x"3b381703", 
    x"3b389bc3", 
    x"3b392144", 
    x"3b39a786", 
    x"3b3a2e8c", 
    x"3b3ab656", 
    x"3b3b3ee7", 
    x"3b3bc841", 
    x"3b3c5264", 
    x"3b3cdd53", 
    x"3b3d6910", 
    x"3b3df59d", 
    x"3b3e82fa", 
    x"3b3f112b", 
    x"3b3fa030", 
    x"3b40300c", 
    x"3b40c0c1", 
    x"3b415250", 
    x"3b41e4bc", 
    x"3b427806", 
    x"3b430c31", 
    x"3b43a13e", 
    x"3b443730", 
    x"3b44ce08", 
    x"3b4565c8", 
    x"3b45fe74", 
    x"3b46980c", 
    x"3b473294", 
    x"3b47ce0c", 
    x"3b486a79", 
    x"3b4907da", 
    x"3b49a634", 
    x"3b4a4588", 
    x"3b4ae5d8", 
    x"3b4b8728", 
    x"3b4c2978", 
    x"3b4ccccd", 
    x"3b4d7127", 
    x"3b4e168a", 
    x"3b4ebcf9", 
    x"3b4f6475", 
    x"3b500d01", 
    x"3b50b6a0", 
    x"3b516154", 
    x"3b520d21", 
    x"3b52ba08", 
    x"3b53680d", 
    x"3b541733", 
    x"3b54c77b", 
    x"3b5578e9", 
    x"3b562b81", 
    x"3b56df44", 
    x"3b579436", 
    x"3b584a5a", 
    x"3b5901b2", 
    x"3b59ba42", 
    x"3b5a740e", 
    x"3b5b2f17", 
    x"3b5beb62", 
    x"3b5ca8f1", 
    x"3b5d67c9", 
    x"3b5e27eb", 
    x"3b5ee95c", 
    x"3b5fac1f", 
    x"3b607038", 
    x"3b6135aa", 
    x"3b61fc78", 
    x"3b62c4a7", 
    x"3b638e39", 
    x"3b645933", 
    x"3b652598", 
    x"3b65f36d", 
    x"3b66c2b4", 
    x"3b679373", 
    x"3b6865ac", 
    x"3b693965", 
    x"3b6a0ea1", 
    x"3b6ae564", 
    x"3b6bbdb3", 
    x"3b6c9791", 
    x"3b6d7304", 
    x"3b6e500f", 
    x"3b6f2eb7", 
    x"3b700f01", 
    x"3b70f0f1", 
    x"3b71d48c", 
    x"3b72b9d6", 
    x"3b73a0d5", 
    x"3b74898d", 
    x"3b757404", 
    x"3b76603e", 
    x"3b774e40", 
    x"3b783e10", 
    x"3b792fb2", 
    x"3b7a232d", 
    x"3b7b1885", 
    x"3b7c0fc1", 
    x"3b7d08e5", 
    x"3b7e03f8", 
    x"3b7f00ff", 
    x"3b800000", 
    x"3b808081", 
    x"3b810204", 
    x"3b81848e", 
    x"3b820821", 
    x"3b828cc0", 
    x"3b83126f", 
    x"3b839930", 
    x"3b842108", 
    x"3b84a9fa", 
    x"3b853408", 
    x"3b85bf37", 
    x"3b864b8a", 
    x"3b86d905", 
    x"3b8767ab", 
    x"3b87f781", 
    x"3b888889", 
    x"3b891ac7", 
    x"3b89ae41", 
    x"3b8a42f8", 
    x"3b8ad8f3", 
    x"3b8b7034", 
    x"3b8c08c1", 
    x"3b8ca29c", 
    x"3b8d3dcb", 
    x"3b8dda52", 
    x"3b8e7835", 
    x"3b8f177a", 
    x"3b8fb824", 
    x"3b905a38", 
    x"3b90fdbc", 
    x"3b91a2b4", 
    x"3b924925", 
    x"3b92f114", 
    x"3b939a86", 
    x"3b944581", 
    x"3b94f209", 
    x"3b95a025", 
    x"3b964fda", 
    x"3b97012e", 
    x"3b97b426", 
    x"3b9868c8", 
    x"3b991f1a", 
    x"3b99d723", 
    x"3b9a90e8", 
    x"3b9b4c70", 
    x"3b9c09c1", 
    x"3b9cc8e1", 
    x"3b9d89d9", 
    x"3b9e4cad", 
    x"3b9f1166", 
    x"3b9fd80a", 
    x"3ba0a0a1", 
    x"3ba16b31", 
    x"3ba237c3", 
    x"3ba3065e", 
    x"3ba3d70a", 
    x"3ba4a9cf", 
    x"3ba57eb5", 
    x"3ba655c4", 
    x"3ba72f05", 
    x"3ba80a81", 
    x"3ba8e83f", 
    x"3ba9c84a", 
    x"3baaaaab", 
    x"3bab8f6a", 
    x"3bac7692", 
    x"3bad602b", 
    x"3bae4c41", 
    x"3baf3ade", 
    x"3bb02c0b", 
    x"3bb11fd4", 
    x"3bb21643", 
    x"3bb30f63", 
    x"3bb40b41", 
    x"3bb509e7", 
    x"3bb60b61", 
    x"3bb70fbb", 
    x"3bb81703", 
    x"3bb92144", 
    x"3bba2e8c", 
    x"3bbb3ee7", 
    x"3bbc5264", 
    x"3bbd6910", 
    x"3bbe82fa", 
    x"3bbfa030", 
    x"3bc0c0c1", 
    x"3bc1e4bc", 
    x"3bc30c31", 
    x"3bc43730", 
    x"3bc565c8", 
    x"3bc6980c", 
    x"3bc7ce0c", 
    x"3bc907da", 
    x"3bca4588", 
    x"3bcb8728", 
    x"3bcccccd", 
    x"3bce168a", 
    x"3bcf6475", 
    x"3bd0b6a0", 
    x"3bd20d21", 
    x"3bd3680d", 
    x"3bd4c77b", 
    x"3bd62b81", 
    x"3bd79436", 
    x"3bd901b2", 
    x"3bda740e", 
    x"3bdbeb62", 
    x"3bdd67c9", 
    x"3bdee95c", 
    x"3be07038", 
    x"3be1fc78", 
    x"3be38e39", 
    x"3be52598", 
    x"3be6c2b4", 
    x"3be865ac", 
    x"3bea0ea1", 
    x"3bebbdb3", 
    x"3bed7304", 
    x"3bef2eb7", 
    x"3bf0f0f1", 
    x"3bf2b9d6", 
    x"3bf4898d", 
    x"3bf6603e", 
    x"3bf83e10", 
    x"3bfa232d", 
    x"3bfc0fc1", 
    x"3bfe03f8", 
    x"3c000000", 
    x"3c010204", 
    x"3c020821", 
    x"3c03126f", 
    x"3c042108", 
    x"3c053408", 
    x"3c064b8a", 
    x"3c0767ab", 
    x"3c088889", 
    x"3c09ae41", 
    x"3c0ad8f3", 
    x"3c0c08c1", 
    x"3c0d3dcb", 
    x"3c0e7835", 
    x"3c0fb824", 
    x"3c10fdbc", 
    x"3c124925", 
    x"3c139a86", 
    x"3c14f209", 
    x"3c164fda", 
    x"3c17b426", 
    x"3c191f1a", 
    x"3c1a90e8", 
    x"3c1c09c1", 
    x"3c1d89d9", 
    x"3c1f1166", 
    x"3c20a0a1", 
    x"3c2237c3", 
    x"3c23d70a", 
    x"3c257eb5", 
    x"3c272f05", 
    x"3c28e83f", 
    x"3c2aaaab", 
    x"3c2c7692", 
    x"3c2e4c41", 
    x"3c302c0b", 
    x"3c321643", 
    x"3c340b41", 
    x"3c360b61", 
    x"3c381703", 
    x"3c3a2e8c", 
    x"3c3c5264", 
    x"3c3e82fa", 
    x"3c40c0c1", 
    x"3c430c31", 
    x"3c4565c8", 
    x"3c47ce0c", 
    x"3c4a4588", 
    x"3c4ccccd", 
    x"3c4f6475", 
    x"3c520d21", 
    x"3c54c77b", 
    x"3c579436", 
    x"3c5a740e", 
    x"3c5d67c9", 
    x"3c607038", 
    x"3c638e39", 
    x"3c66c2b4", 
    x"3c6a0ea1", 
    x"3c6d7304", 
    x"3c70f0f1", 
    x"3c74898d", 
    x"3c783e10", 
    x"3c7c0fc1", 
    x"3c800000", 
    x"3c820821", 
    x"3c842108", 
    x"3c864b8a", 
    x"3c888889", 
    x"3c8ad8f3", 
    x"3c8d3dcb", 
    x"3c8fb824", 
    x"3c924925", 
    x"3c94f209", 
    x"3c97b426", 
    x"3c9a90e8", 
    x"3c9d89d9", 
    x"3ca0a0a1", 
    x"3ca3d70a", 
    x"3ca72f05", 
    x"3caaaaab", 
    x"3cae4c41", 
    x"3cb21643", 
    x"3cb60b61", 
    x"3cba2e8c", 
    x"3cbe82fa", 
    x"3cc30c31", 
    x"3cc7ce0c", 
    x"3ccccccd", 
    x"3cd20d21", 
    x"3cd79436", 
    x"3cdd67c9", 
    x"3ce38e39", 
    x"3cea0ea1", 
    x"3cf0f0f1", 
    x"3cf83e10", 
    x"3d000000", 
    x"3d042108", 
    x"3d088889", 
    x"3d0d3dcb", 
    x"3d124925", 
    x"3d17b426", 
    x"3d1d89d9", 
    x"3d23d70a", 
    x"3d2aaaab", 
    x"3d321643", 
    x"3d3a2e8c", 
    x"3d430c31", 
    x"3d4ccccd", 
    x"3d579436", 
    x"3d638e39", 
    x"3d70f0f1", 
    x"3d800000", 
    x"3d888889", 
    x"3d924925", 
    x"3d9d89d9", 
    x"3daaaaab", 
    x"3dba2e8c", 
    x"3dcccccd", 
    x"3de38e39", 
    x"3e000000", 
    x"3e124925", 
    x"3e2aaaab", 
    x"3e4ccccd", 
    x"3e800000", 
    x"3eaaaaab", 
    x"3f000000", 
    x"3f800000", 
    x"00000000"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
