-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom3 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom3; 
 
architecture behavioral of inv_rom3 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"3a2aaaab", 
    x"3a2a8e3e", 
    x"3a2a71da", 
    x"3a2a5580", 
    x"3a2a392f", 
    x"3a2a1ce8", 
    x"3a2a00aa", 
    x"3a29e475", 
    x"3a29c84a", 
    x"3a29ac28", 
    x"3a299010", 
    x"3a297401", 
    x"3a2957fb", 
    x"3a293bfe", 
    x"3a29200b", 
    x"3a290420", 
    x"3a28e83f", 
    x"3a28cc68", 
    x"3a28b099", 
    x"3a2894d3", 
    x"3a287917", 
    x"3a285d64", 
    x"3a2841ba", 
    x"3a282619", 
    x"3a280a81", 
    x"3a27eef2", 
    x"3a27d36c", 
    x"3a27b7ef", 
    x"3a279c7b", 
    x"3a278110", 
    x"3a2765ae", 
    x"3a274a55", 
    x"3a272f05", 
    x"3a2713be", 
    x"3a26f880", 
    x"3a26dd4a", 
    x"3a26c21e", 
    x"3a26a6fa", 
    x"3a268bdf", 
    x"3a2670cd", 
    x"3a2655c4", 
    x"3a263ac4", 
    x"3a261fcc", 
    x"3a2604dd", 
    x"3a25e9f7", 
    x"3a25cf19", 
    x"3a25b445", 
    x"3a259978", 
    x"3a257eb5", 
    x"3a2563fa", 
    x"3a254948", 
    x"3a252e9e", 
    x"3a2513fd", 
    x"3a24f965", 
    x"3a24ded5", 
    x"3a24c44e", 
    x"3a24a9cf", 
    x"3a248f59", 
    x"3a2474eb", 
    x"3a245a86", 
    x"3a244029", 
    x"3a2425d5", 
    x"3a240b89", 
    x"3a23f145", 
    x"3a23d70a", 
    x"3a23bcd8", 
    x"3a23a2ad", 
    x"3a23888b", 
    x"3a236e72", 
    x"3a235460", 
    x"3a233a57", 
    x"3a232057", 
    x"3a23065e", 
    x"3a22ec6e", 
    x"3a22d286", 
    x"3a22b8a7", 
    x"3a229ecf", 
    x"3a228500", 
    x"3a226b39", 
    x"3a22517a", 
    x"3a2237c3", 
    x"3a221e15", 
    x"3a22046e", 
    x"3a21ead0", 
    x"3a21d13a", 
    x"3a21b7ab", 
    x"3a219e25", 
    x"3a2184a7", 
    x"3a216b31", 
    x"3a2151c3", 
    x"3a21385d", 
    x"3a211eff", 
    x"3a2105a9", 
    x"3a20ec5b", 
    x"3a20d315", 
    x"3a20b9d7", 
    x"3a20a0a1", 
    x"3a208772", 
    x"3a206e4c", 
    x"3a20552d", 
    x"3a203c17", 
    x"3a202308", 
    x"3a200a01", 
    x"3a1ff101", 
    x"3a1fd80a", 
    x"3a1fbf1a", 
    x"3a1fa633", 
    x"3a1f8d52", 
    x"3a1f747a", 
    x"3a1f5ba9", 
    x"3a1f42e1", 
    x"3a1f2a1f", 
    x"3a1f1166", 
    x"3a1ef8b4", 
    x"3a1ee00a", 
    x"3a1ec767", 
    x"3a1eaecd", 
    x"3a1e9639", 
    x"3a1e7dae", 
    x"3a1e652a", 
    x"3a1e4cad", 
    x"3a1e3438", 
    x"3a1e1bcb", 
    x"3a1e0365", 
    x"3a1deb07", 
    x"3a1dd2b0", 
    x"3a1dba61", 
    x"3a1da219", 
    x"3a1d89d9", 
    x"3a1d71a0", 
    x"3a1d596e", 
    x"3a1d4144", 
    x"3a1d2922", 
    x"3a1d1107", 
    x"3a1cf8f3", 
    x"3a1ce0e6", 
    x"3a1cc8e1", 
    x"3a1cb0e4", 
    x"3a1c98ed", 
    x"3a1c80fe", 
    x"3a1c6917", 
    x"3a1c5136", 
    x"3a1c395d", 
    x"3a1c218b", 
    x"3a1c09c1", 
    x"3a1bf1fd", 
    x"3a1bda41", 
    x"3a1bc28c", 
    x"3a1baadf", 
    x"3a1b9338", 
    x"3a1b7b99", 
    x"3a1b6401", 
    x"3a1b4c70", 
    x"3a1b34e6", 
    x"3a1b1d63", 
    x"3a1b05e7", 
    x"3a1aee73", 
    x"3a1ad706", 
    x"3a1abf9f", 
    x"3a1aa840", 
    x"3a1a90e8", 
    x"3a1a7997", 
    x"3a1a624d", 
    x"3a1a4b09", 
    x"3a1a33cd", 
    x"3a1a1c98", 
    x"3a1a056a", 
    x"3a19ee43", 
    x"3a19d723", 
    x"3a19c00a", 
    x"3a19a8f7", 
    x"3a1991ec", 
    x"3a197ae7", 
    x"3a1963ea", 
    x"3a194cf3", 
    x"3a193603", 
    x"3a191f1a", 
    x"3a190838", 
    x"3a18f15d", 
    x"3a18da88", 
    x"3a18c3bb", 
    x"3a18acf4", 
    x"3a189634", 
    x"3a187f7b", 
    x"3a1868c8", 
    x"3a18521c", 
    x"3a183b77", 
    x"3a1824d9", 
    x"3a180e41", 
    x"3a17f7b0", 
    x"3a17e126", 
    x"3a17caa3", 
    x"3a17b426", 
    x"3a179db0", 
    x"3a178740", 
    x"3a1770d7", 
    x"3a175a75", 
    x"3a174419", 
    x"3a172dc4", 
    x"3a171776", 
    x"3a17012e", 
    x"3a16eaed", 
    x"3a16d4b2", 
    x"3a16be7e", 
    x"3a16a850", 
    x"3a169229", 
    x"3a167c08", 
    x"3a1665ee", 
    x"3a164fda", 
    x"3a1639cd", 
    x"3a1623c7", 
    x"3a160dc6", 
    x"3a15f7cc", 
    x"3a15e1d9", 
    x"3a15cbec", 
    x"3a15b606", 
    x"3a15a025", 
    x"3a158a4c", 
    x"3a157478", 
    x"3a155eab", 
    x"3a1548e5", 
    x"3a153324", 
    x"3a151d6a", 
    x"3a1507b7", 
    x"3a14f209", 
    x"3a14dc62", 
    x"3a14c6c2", 
    x"3a14b127", 
    x"3a149b93", 
    x"3a148605", 
    x"3a14707d", 
    x"3a145afc", 
    x"3a144581", 
    x"3a14300c", 
    x"3a141a9d", 
    x"3a140534", 
    x"3a13efd2", 
    x"3a13da76", 
    x"3a13c51f", 
    x"3a13afd0", 
    x"3a139a86", 
    x"3a138542", 
    x"3a137005", 
    x"3a135acd", 
    x"3a13459c", 
    x"3a133071", 
    x"3a131b4c", 
    x"3a13062d", 
    x"3a12f114", 
    x"3a12dc01", 
    x"3a12c6f4", 
    x"3a12b1ed", 
    x"3a129cec", 
    x"3a1287f1", 
    x"3a1272fc", 
    x"3a125e0d", 
    x"3a124925", 
    x"3a123442", 
    x"3a121f65", 
    x"3a120a8e", 
    x"3a11f5bd", 
    x"3a11e0f2", 
    x"3a11cc2c", 
    x"3a11b76d", 
    x"3a11a2b4", 
    x"3a118e00", 
    x"3a117953", 
    x"3a1164ab", 
    x"3a115009", 
    x"3a113b6d", 
    x"3a1126d7", 
    x"3a111247", 
    x"3a10fdbc", 
    x"3a10e937", 
    x"3a10d4b8", 
    x"3a10c03f", 
    x"3a10abcc", 
    x"3a10975e", 
    x"3a1082f7", 
    x"3a106e95", 
    x"3a105a38", 
    x"3a1045e2", 
    x"3a103191", 
    x"3a101d46", 
    x"3a100901", 
    x"3a0ff4c1", 
    x"3a0fe087", 
    x"3a0fcc53", 
    x"3a0fb824", 
    x"3a0fa3fb", 
    x"3a0f8fd8", 
    x"3a0f7bba", 
    x"3a0f67a2", 
    x"3a0f538f", 
    x"3a0f3f83", 
    x"3a0f2b7b", 
    x"3a0f177a", 
    x"3a0f037e", 
    x"3a0eef87", 
    x"3a0edb97", 
    x"3a0ec7ab", 
    x"3a0eb3c5", 
    x"3a0e9fe5", 
    x"3a0e8c0b", 
    x"3a0e7835", 
    x"3a0e6466", 
    x"3a0e509c", 
    x"3a0e3cd7", 
    x"3a0e2918", 
    x"3a0e155e", 
    x"3a0e01aa", 
    x"3a0dedfb", 
    x"3a0dda52", 
    x"3a0dc6ae", 
    x"3a0db310", 
    x"3a0d9f77", 
    x"3a0d8be3", 
    x"3a0d7855", 
    x"3a0d64cc", 
    x"3a0d5149", 
    x"3a0d3dcb", 
    x"3a0d2a52", 
    x"3a0d16df", 
    x"3a0d0371", 
    x"3a0cf009", 
    x"3a0cdca6", 
    x"3a0cc948", 
    x"3a0cb5ef", 
    x"3a0ca29c", 
    x"3a0c8f4e", 
    x"3a0c7c05", 
    x"3a0c68c2", 
    x"3a0c5584", 
    x"3a0c424b", 
    x"3a0c2f18", 
    x"3a0c1bea", 
    x"3a0c08c1", 
    x"3a0bf59d", 
    x"3a0be27e", 
    x"3a0bcf65", 
    x"3a0bbc51", 
    x"3a0ba942", 
    x"3a0b9638", 
    x"3a0b8334", 
    x"3a0b7034", 
    x"3a0b5d3a", 
    x"3a0b4a45", 
    x"3a0b3755", 
    x"3a0b246b", 
    x"3a0b1185", 
    x"3a0afea5", 
    x"3a0aebc9", 
    x"3a0ad8f3", 
    x"3a0ac622", 
    x"3a0ab356", 
    x"3a0aa08f", 
    x"3a0a8dcd", 
    x"3a0a7b10", 
    x"3a0a6859", 
    x"3a0a55a6", 
    x"3a0a42f8", 
    x"3a0a3050", 
    x"3a0a1dac", 
    x"3a0a0b0e", 
    x"3a09f874", 
    x"3a09e5e0", 
    x"3a09d350", 
    x"3a09c0c6", 
    x"3a09ae41", 
    x"3a099bc0", 
    x"3a098944", 
    x"3a0976ce", 
    x"3a09645c", 
    x"3a0951f0", 
    x"3a093f88", 
    x"3a092d25", 
    x"3a091ac7", 
    x"3a09086e", 
    x"3a08f61a", 
    x"3a08e3cb", 
    x"3a08d181", 
    x"3a08bf3b", 
    x"3a08acfb", 
    x"3a089abf", 
    x"3a088889", 
    x"3a087657", 
    x"3a08642a", 
    x"3a085201", 
    x"3a083fde", 
    x"3a082dbf", 
    x"3a081ba6", 
    x"3a080991", 
    x"3a07f781", 
    x"3a07e575", 
    x"3a07d36f", 
    x"3a07c16d", 
    x"3a07af70", 
    x"3a079d78", 
    x"3a078b84", 
    x"3a077995", 
    x"3a0767ab", 
    x"3a0755c6", 
    x"3a0743e6", 
    x"3a07320a", 
    x"3a072033", 
    x"3a070e60", 
    x"3a06fc93", 
    x"3a06eaca", 
    x"3a06d905", 
    x"3a06c746", 
    x"3a06b58b", 
    x"3a06a3d4", 
    x"3a069223", 
    x"3a068076", 
    x"3a066ecd", 
    x"3a065d2a", 
    x"3a064b8a", 
    x"3a0639f0", 
    x"3a06285a", 
    x"3a0616c9", 
    x"3a06053c", 
    x"3a05f3b4", 
    x"3a05e231", 
    x"3a05d0b2", 
    x"3a05bf37", 
    x"3a05adc2", 
    x"3a059c50", 
    x"3a058ae4", 
    x"3a05797c", 
    x"3a056818", 
    x"3a0556b9", 
    x"3a05455e", 
    x"3a053408", 
    x"3a0522b7", 
    x"3a05116a", 
    x"3a050021", 
    x"3a04eedd", 
    x"3a04dd9e", 
    x"3a04cc63", 
    x"3a04bb2c", 
    x"3a04a9fa", 
    x"3a0498cc", 
    x"3a0487a3", 
    x"3a04767e", 
    x"3a04655e", 
    x"3a045442", 
    x"3a04432a", 
    x"3a043217", 
    x"3a042108", 
    x"3a040ffe", 
    x"3a03fef8", 
    x"3a03edf6", 
    x"3a03dcf9", 
    x"3a03cc01", 
    x"3a03bb0c", 
    x"3a03aa1c", 
    x"3a039930", 
    x"3a038849", 
    x"3a037766", 
    x"3a036687", 
    x"3a0355ad", 
    x"3a0344d7", 
    x"3a033405", 
    x"3a032338", 
    x"3a03126f", 
    x"3a0301aa", 
    x"3a02f0e9", 
    x"3a02e02d", 
    x"3a02cf75", 
    x"3a02bec1", 
    x"3a02ae12", 
    x"3a029d67", 
    x"3a028cc0", 
    x"3a027c1d", 
    x"3a026b7f", 
    x"3a025ae4", 
    x"3a024a4e", 
    x"3a0239bd", 
    x"3a02292f", 
    x"3a0218a6", 
    x"3a020821", 
    x"3a01f7a0", 
    x"3a01e723", 
    x"3a01d6aa", 
    x"3a01c636", 
    x"3a01b5c5", 
    x"3a01a559", 
    x"3a0194f1", 
    x"3a01848e", 
    x"3a01742e", 
    x"3a0163d3", 
    x"3a01537b", 
    x"3a014328", 
    x"3a0132d9", 
    x"3a01228e", 
    x"3a011247", 
    x"3a010204", 
    x"3a00f1c5", 
    x"3a00e18b", 
    x"3a00d154", 
    x"3a00c122", 
    x"3a00b0f3", 
    x"3a00a0c9", 
    x"3a0090a3", 
    x"3a008081", 
    x"3a007062", 
    x"3a006048", 
    x"3a005032", 
    x"3a004020", 
    x"3a003012", 
    x"3a002008", 
    x"3a001002"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
