-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom8 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom8; 
 
architecture behavioral of inv_rom8 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"39800000", 
    x"397ff001", 
    x"397fe004", 
    x"397fd009", 
    x"397fc010", 
    x"397fb019", 
    x"397fa024", 
    x"397f9031", 
    x"397f8040", 
    x"397f7051", 
    x"397f6064", 
    x"397f5079", 
    x"397f4090", 
    x"397f30a8", 
    x"397f20c3", 
    x"397f10e0", 
    x"397f00ff", 
    x"397ef120", 
    x"397ee143", 
    x"397ed167", 
    x"397ec18e", 
    x"397eb1b7", 
    x"397ea1e1", 
    x"397e920e", 
    x"397e823d", 
    x"397e726d", 
    x"397e62a0", 
    x"397e52d4", 
    x"397e430b", 
    x"397e3343", 
    x"397e237d", 
    x"397e13ba", 
    x"397e03f8", 
    x"397df438", 
    x"397de47a", 
    x"397dd4bf", 
    x"397dc505", 
    x"397db54d", 
    x"397da597", 
    x"397d95e3", 
    x"397d8631", 
    x"397d7680", 
    x"397d66d2", 
    x"397d5726", 
    x"397d477b", 
    x"397d37d3", 
    x"397d282d", 
    x"397d1888", 
    x"397d08e5", 
    x"397cf945", 
    x"397ce9a6", 
    x"397cda09", 
    x"397cca6e", 
    x"397cbad5", 
    x"397cab3e", 
    x"397c9ba9", 
    x"397c8c16", 
    x"397c7c84", 
    x"397c6cf5", 
    x"397c5d68", 
    x"397c4ddc", 
    x"397c3e52", 
    x"397c2ecb", 
    x"397c1f45", 
    x"397c0fc1", 
    x"397c003f", 
    x"397bf0bf", 
    x"397be141", 
    x"397bd1c4", 
    x"397bc24a", 
    x"397bb2d2", 
    x"397ba35b", 
    x"397b93e6", 
    x"397b8474", 
    x"397b7503", 
    x"397b6594", 
    x"397b5627", 
    x"397b46bc", 
    x"397b3752", 
    x"397b27eb", 
    x"397b1885", 
    x"397b0922", 
    x"397af9c0", 
    x"397aea60", 
    x"397adb02", 
    x"397acba6", 
    x"397abc4c", 
    x"397aacf4", 
    x"397a9d9d", 
    x"397a8e49", 
    x"397a7ef6", 
    x"397a6fa5", 
    x"397a6056", 
    x"397a5109", 
    x"397a41be", 
    x"397a3274", 
    x"397a232d", 
    x"397a13e7", 
    x"397a04a4", 
    x"3979f562", 
    x"3979e622", 
    x"3979d6e4", 
    x"3979c7a7", 
    x"3979b86d", 
    x"3979a934", 
    x"397999fd", 
    x"39798ac9", 
    x"39797b96", 
    x"39796c64", 
    x"39795d35", 
    x"39794e08", 
    x"39793edc", 
    x"39792fb2", 
    x"3979208a", 
    x"39791164", 
    x"39790240", 
    x"3978f31d", 
    x"3978e3fd", 
    x"3978d4de", 
    x"3978c5c1", 
    x"3978b6a6", 
    x"3978a78d", 
    x"39789876", 
    x"39788960", 
    x"39787a4c", 
    x"39786b3a", 
    x"39785c2a", 
    x"39784d1c", 
    x"39783e10", 
    x"39782f05", 
    x"39781ffc", 
    x"397810f5", 
    x"397801f0", 
    x"3977f2ed", 
    x"3977e3eb", 
    x"3977d4eb", 
    x"3977c5ee", 
    x"3977b6f2", 
    x"3977a7f7", 
    x"397798ff", 
    x"39778a08", 
    x"39777b13", 
    x"39776c20", 
    x"39775d2f", 
    x"39774e40", 
    x"39773f52", 
    x"39773066", 
    x"3977217c", 
    x"39771294", 
    x"397703ae", 
    x"3976f4c9", 
    x"3976e5e6", 
    x"3976d705", 
    x"3976c826", 
    x"3976b949", 
    x"3976aa6d", 
    x"39769b93", 
    x"39768cbb", 
    x"39767de5", 
    x"39766f10", 
    x"3976603e", 
    x"3976516d", 
    x"3976429e", 
    x"397633d0", 
    x"39762505", 
    x"3976163b", 
    x"39760773", 
    x"3975f8ac", 
    x"3975e9e8", 
    x"3975db25", 
    x"3975cc64", 
    x"3975bda5", 
    x"3975aee8", 
    x"3975a02c", 
    x"39759172", 
    x"397582ba", 
    x"39757404", 
    x"3975654f", 
    x"3975569c", 
    x"397547eb", 
    x"3975393c", 
    x"39752a8f", 
    x"39751be3", 
    x"39750d39", 
    x"3974fe91", 
    x"3974efea", 
    x"3974e145", 
    x"3974d2a2", 
    x"3974c401", 
    x"3974b561", 
    x"3974a6c4", 
    x"39749828", 
    x"3974898d", 
    x"39747af5", 
    x"39746c5e", 
    x"39745dc9", 
    x"39744f36", 
    x"397440a4", 
    x"39743214", 
    x"39742386", 
    x"397414fa", 
    x"3974066f", 
    x"3973f7e6", 
    x"3973e95f", 
    x"3973dada", 
    x"3973cc56", 
    x"3973bdd4", 
    x"3973af54", 
    x"3973a0d5", 
    x"39739258", 
    x"397383dd", 
    x"39737564", 
    x"397366ec", 
    x"39735876", 
    x"39734a02", 
    x"39733b90", 
    x"39732d1f", 
    x"39731eb0", 
    x"39731042", 
    x"397301d7", 
    x"3972f36d", 
    x"3972e505", 
    x"3972d69e", 
    x"3972c839", 
    x"3972b9d6", 
    x"3972ab75", 
    x"39729d15", 
    x"39728eb7", 
    x"3972805b", 
    x"39727200", 
    x"397263a7", 
    x"39725550", 
    x"397246fb", 
    x"397238a7", 
    x"39722a55", 
    x"39721c04", 
    x"39720db6", 
    x"3971ff69", 
    x"3971f11d", 
    x"3971e2d4", 
    x"3971d48c", 
    x"3971c646", 
    x"3971b801", 
    x"3971a9be", 
    x"39719b7d", 
    x"39718d3d", 
    x"39717eff", 
    x"397170c3", 
    x"39716289", 
    x"39715450", 
    x"39714619", 
    x"397137e3", 
    x"397129af", 
    x"39711b7d", 
    x"39710d4d", 
    x"3970ff1e", 
    x"3970f0f1", 
    x"3970e2c5", 
    x"3970d49c", 
    x"3970c674", 
    x"3970b84d", 
    x"3970aa28", 
    x"39709c05", 
    x"39708de4", 
    x"39707fc4", 
    x"397071a6", 
    x"39706389", 
    x"3970556e", 
    x"39704755", 
    x"3970393e", 
    x"39702b28", 
    x"39701d14", 
    x"39700f01", 
    x"397000f0", 
    x"396ff2e1", 
    x"396fe4d3", 
    x"396fd6c7", 
    x"396fc8bd", 
    x"396fbab4", 
    x"396facad", 
    x"396f9ea8", 
    x"396f90a4", 
    x"396f82a2", 
    x"396f74a1", 
    x"396f66a2", 
    x"396f58a5", 
    x"396f4aa9", 
    x"396f3caf", 
    x"396f2eb7", 
    x"396f20c0", 
    x"396f12cb", 
    x"396f04d8", 
    x"396ef6e6", 
    x"396ee8f6", 
    x"396edb07", 
    x"396ecd1a", 
    x"396ebf2f", 
    x"396eb145", 
    x"396ea35d", 
    x"396e9577", 
    x"396e8792", 
    x"396e79af", 
    x"396e6bcd", 
    x"396e5ded", 
    x"396e500f", 
    x"396e4232", 
    x"396e3457", 
    x"396e267d", 
    x"396e18a6", 
    x"396e0acf", 
    x"396dfcfb", 
    x"396def27", 
    x"396de156", 
    x"396dd386", 
    x"396dc5b8", 
    x"396db7eb", 
    x"396daa20", 
    x"396d9c57", 
    x"396d8e8f", 
    x"396d80c8", 
    x"396d7304", 
    x"396d6541", 
    x"396d577f", 
    x"396d49bf", 
    x"396d3c01", 
    x"396d2e44", 
    x"396d2089", 
    x"396d12d0", 
    x"396d0518", 
    x"396cf761", 
    x"396ce9ac", 
    x"396cdbf9", 
    x"396cce48", 
    x"396cc098", 
    x"396cb2e9", 
    x"396ca53c", 
    x"396c9791", 
    x"396c89e7", 
    x"396c7c3f", 
    x"396c6e99", 
    x"396c60f4", 
    x"396c5350", 
    x"396c45af", 
    x"396c380e", 
    x"396c2a70", 
    x"396c1cd3", 
    x"396c0f37", 
    x"396c019d", 
    x"396bf405", 
    x"396be66e", 
    x"396bd8d9", 
    x"396bcb45", 
    x"396bbdb3", 
    x"396bb022", 
    x"396ba293", 
    x"396b9506", 
    x"396b877a", 
    x"396b79ef", 
    x"396b6c67", 
    x"396b5edf", 
    x"396b515a", 
    x"396b43d5", 
    x"396b3653", 
    x"396b28d2", 
    x"396b1b52", 
    x"396b0dd5", 
    x"396b0058", 
    x"396af2dd", 
    x"396ae564", 
    x"396ad7ec", 
    x"396aca76", 
    x"396abd01", 
    x"396aaf8e", 
    x"396aa21d", 
    x"396a94ad", 
    x"396a873e", 
    x"396a79d1", 
    x"396a6c66", 
    x"396a5efc", 
    x"396a5194", 
    x"396a442d", 
    x"396a36c8", 
    x"396a2964", 
    x"396a1c02", 
    x"396a0ea1", 
    x"396a0142", 
    x"3969f3e4", 
    x"3969e688", 
    x"3969d92d", 
    x"3969cbd4", 
    x"3969be7d", 
    x"3969b127", 
    x"3969a3d2", 
    x"3969967f", 
    x"3969892e", 
    x"39697bde", 
    x"39696e90", 
    x"39696143", 
    x"396953f7", 
    x"396946ad", 
    x"39693965", 
    x"39692c1e", 
    x"39691ed9", 
    x"39691195", 
    x"39690453", 
    x"3968f712", 
    x"3968e9d3", 
    x"3968dc95", 
    x"3968cf59", 
    x"3968c21e", 
    x"3968b4e5", 
    x"3968a7ad", 
    x"39689a77", 
    x"39688d42", 
    x"3968800f", 
    x"396872dd", 
    x"396865ac", 
    x"3968587e", 
    x"39684b50", 
    x"39683e25", 
    x"396830fa", 
    x"396823d2", 
    x"396816aa", 
    x"39680984", 
    x"3967fc60", 
    x"3967ef3d", 
    x"3967e21c", 
    x"3967d4fc", 
    x"3967c7de", 
    x"3967bac1", 
    x"3967ada5", 
    x"3967a08b", 
    x"39679373", 
    x"3967865c", 
    x"39677946", 
    x"39676c32", 
    x"39675f20", 
    x"3967520f", 
    x"396744ff", 
    x"396737f1", 
    x"39672ae4", 
    x"39671dd9", 
    x"396710d0", 
    x"396703c7", 
    x"3966f6c1", 
    x"3966e9bb", 
    x"3966dcb8", 
    x"3966cfb5", 
    x"3966c2b4", 
    x"3966b5b5", 
    x"3966a8b7", 
    x"39669bba", 
    x"39668ebf", 
    x"396681c6", 
    x"396674ce", 
    x"396667d7", 
    x"39665ae2", 
    x"39664dee", 
    x"396640fc", 
    x"3966340b", 
    x"3966271c", 
    x"39661a2e", 
    x"39660d41", 
    x"39660056", 
    x"3965f36d", 
    x"3965e685", 
    x"3965d99e", 
    x"3965ccb9", 
    x"3965bfd5", 
    x"3965b2f3", 
    x"3965a612", 
    x"39659932", 
    x"39658c54", 
    x"39657f78", 
    x"3965729d", 
    x"396565c3", 
    x"396558eb", 
    x"39654c14", 
    x"39653f3f", 
    x"3965326b", 
    x"39652598", 
    x"396518c7", 
    x"39650bf8", 
    x"3964ff29", 
    x"3964f25d", 
    x"3964e591", 
    x"3964d8c7", 
    x"3964cbff", 
    x"3964bf38", 
    x"3964b272", 
    x"3964a5ae", 
    x"396498eb", 
    x"39648c2a", 
    x"39647f6a", 
    x"396472ac", 
    x"396465ee", 
    x"39645933", 
    x"39644c79", 
    x"39643fc0", 
    x"39643308", 
    x"39642652", 
    x"3964199e", 
    x"39640ceb", 
    x"39640039", 
    x"3963f389", 
    x"3963e6da", 
    x"3963da2c", 
    x"3963cd80", 
    x"3963c0d6", 
    x"3963b42c", 
    x"3963a784", 
    x"39639ade"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
