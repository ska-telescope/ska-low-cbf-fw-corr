-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom6 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom6; 
 
architecture behavioral of inv_rom6 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"39925398", 
    x"39925e0d", 
    x"39926884", 
    x"399272fc", 
    x"39927d76", 
    x"399287f1", 
    x"3992926e", 
    x"39929cec", 
    x"3992a76c", 
    x"3992b1ed", 
    x"3992bc6f", 
    x"3992c6f4", 
    x"3992d179", 
    x"3992dc01", 
    x"3992e689", 
    x"3992f114", 
    x"3992fb9f", 
    x"3993062d", 
    x"399310bb", 
    x"39931b4c", 
    x"399325dd", 
    x"39933071", 
    x"39933b06", 
    x"3993459c", 
    x"39935034", 
    x"39935acd", 
    x"39936568", 
    x"39937005", 
    x"39937aa3", 
    x"39938542", 
    x"39938fe3", 
    x"39939a86", 
    x"3993a52a", 
    x"3993afd0", 
    x"3993ba77", 
    x"3993c51f", 
    x"3993cfca", 
    x"3993da76", 
    x"3993e523", 
    x"3993efd2", 
    x"3993fa82", 
    x"39940534", 
    x"39940fe8", 
    x"39941a9d", 
    x"39942553", 
    x"3994300c", 
    x"39943ac5", 
    x"39944581", 
    x"3994503d", 
    x"39945afc", 
    x"399465bc", 
    x"3994707d", 
    x"39947b40", 
    x"39948605", 
    x"399490cb", 
    x"39949b93", 
    x"3994a65c", 
    x"3994b127", 
    x"3994bbf4", 
    x"3994c6c2", 
    x"3994d191", 
    x"3994dc62", 
    x"3994e735", 
    x"3994f209", 
    x"3994fcdf", 
    x"399507b7", 
    x"39951290", 
    x"39951d6a", 
    x"39952847", 
    x"39953324", 
    x"39953e04", 
    x"399548e5", 
    x"399553c7", 
    x"39955eab", 
    x"39956991", 
    x"39957478", 
    x"39957f61", 
    x"39958a4c", 
    x"39959538", 
    x"3995a025", 
    x"3995ab15", 
    x"3995b606", 
    x"3995c0f8", 
    x"3995cbec", 
    x"3995d6e2", 
    x"3995e1d9", 
    x"3995ecd2", 
    x"3995f7cc", 
    x"399602c9", 
    x"39960dc6", 
    x"399618c6", 
    x"399623c7", 
    x"39962ec9", 
    x"399639cd", 
    x"399644d3", 
    x"39964fda", 
    x"39965ae3", 
    x"399665ee", 
    x"399670fa", 
    x"39967c08", 
    x"39968718", 
    x"39969229", 
    x"39969d3c", 
    x"3996a850", 
    x"3996b366", 
    x"3996be7e", 
    x"3996c997", 
    x"3996d4b2", 
    x"3996dfce", 
    x"3996eaed", 
    x"3996f60d", 
    x"3997012e", 
    x"39970c51", 
    x"39971776", 
    x"3997229c", 
    x"39972dc4", 
    x"399738ee", 
    x"39974419", 
    x"39974f46", 
    x"39975a75", 
    x"399765a5", 
    x"399770d7", 
    x"39977c0b", 
    x"39978740", 
    x"39979277", 
    x"39979db0", 
    x"3997a8ea", 
    x"3997b426", 
    x"3997bf64", 
    x"3997caa3", 
    x"3997d5e4", 
    x"3997e126", 
    x"3997ec6b", 
    x"3997f7b0", 
    x"399802f8", 
    x"39980e41", 
    x"3998198c", 
    x"399824d9", 
    x"39983027", 
    x"39983b77", 
    x"399846c9", 
    x"3998521c", 
    x"39985d71", 
    x"399868c8", 
    x"39987420", 
    x"39987f7b", 
    x"39988ad6", 
    x"39989634", 
    x"3998a193", 
    x"3998acf4", 
    x"3998b857", 
    x"3998c3bb", 
    x"3998cf21", 
    x"3998da88", 
    x"3998e5f2", 
    x"3998f15d", 
    x"3998fcca", 
    x"39990838", 
    x"399913a8", 
    x"39991f1a", 
    x"39992a8e", 
    x"39993603", 
    x"3999417a", 
    x"39994cf3", 
    x"3999586e", 
    x"399963ea", 
    x"39996f68", 
    x"39997ae7", 
    x"39998669", 
    x"399991ec", 
    x"39999d71", 
    x"3999a8f7", 
    x"3999b480", 
    x"3999c00a", 
    x"3999cb95", 
    x"3999d723", 
    x"3999e2b2", 
    x"3999ee43", 
    x"3999f9d6", 
    x"399a056a", 
    x"399a1100", 
    x"399a1c98", 
    x"399a2832", 
    x"399a33cd", 
    x"399a3f6b", 
    x"399a4b09", 
    x"399a56aa", 
    x"399a624d", 
    x"399a6df1", 
    x"399a7997", 
    x"399a853e", 
    x"399a90e8", 
    x"399a9c93", 
    x"399aa840", 
    x"399ab3ef", 
    x"399abf9f", 
    x"399acb52", 
    x"399ad706", 
    x"399ae2bb", 
    x"399aee73", 
    x"399afa2c", 
    x"399b05e7", 
    x"399b11a4", 
    x"399b1d63", 
    x"399b2924", 
    x"399b34e6", 
    x"399b40aa", 
    x"399b4c70", 
    x"399b5837", 
    x"399b6401", 
    x"399b6fcc", 
    x"399b7b99", 
    x"399b8768", 
    x"399b9338", 
    x"399b9f0a", 
    x"399baadf", 
    x"399bb6b5", 
    x"399bc28c", 
    x"399bce66", 
    x"399bda41", 
    x"399be61e", 
    x"399bf1fd", 
    x"399bfdde", 
    x"399c09c1", 
    x"399c15a5", 
    x"399c218b", 
    x"399c2d73", 
    x"399c395d", 
    x"399c4549", 
    x"399c5136", 
    x"399c5d25", 
    x"399c6917", 
    x"399c750a", 
    x"399c80fe", 
    x"399c8cf5", 
    x"399c98ed", 
    x"399ca4e8", 
    x"399cb0e4", 
    x"399cbce2", 
    x"399cc8e1", 
    x"399cd4e3", 
    x"399ce0e6", 
    x"399cecec", 
    x"399cf8f3", 
    x"399d04fc", 
    x"399d1107", 
    x"399d1d13", 
    x"399d2922", 
    x"399d3532", 
    x"399d4144", 
    x"399d4d58", 
    x"399d596e", 
    x"399d6586", 
    x"399d71a0", 
    x"399d7dbb", 
    x"399d89d9", 
    x"399d95f8", 
    x"399da219", 
    x"399dae3c", 
    x"399dba61", 
    x"399dc687", 
    x"399dd2b0", 
    x"399ddeda", 
    x"399deb07", 
    x"399df735", 
    x"399e0365", 
    x"399e0f97", 
    x"399e1bcb", 
    x"399e2801", 
    x"399e3438", 
    x"399e4072", 
    x"399e4cad", 
    x"399e58ea", 
    x"399e652a", 
    x"399e716b", 
    x"399e7dae", 
    x"399e89f3", 
    x"399e9639", 
    x"399ea282", 
    x"399eaecd", 
    x"399ebb19", 
    x"399ec767", 
    x"399ed3b8", 
    x"399ee00a", 
    x"399eec5e", 
    x"399ef8b4", 
    x"399f050c", 
    x"399f1166", 
    x"399f1dc2", 
    x"399f2a1f", 
    x"399f367f", 
    x"399f42e1", 
    x"399f4f44", 
    x"399f5ba9", 
    x"399f6811", 
    x"399f747a", 
    x"399f80e5", 
    x"399f8d52", 
    x"399f99c2", 
    x"399fa633", 
    x"399fb2a5", 
    x"399fbf1a", 
    x"399fcb91", 
    x"399fd80a", 
    x"399fe485", 
    x"399ff101", 
    x"399ffd80", 
    x"39a00a01", 
    x"39a01683", 
    x"39a02308", 
    x"39a02f8e", 
    x"39a03c17", 
    x"39a048a1", 
    x"39a0552d", 
    x"39a061bc", 
    x"39a06e4c", 
    x"39a07ade", 
    x"39a08772", 
    x"39a09408", 
    x"39a0a0a1", 
    x"39a0ad3b", 
    x"39a0b9d7", 
    x"39a0c675", 
    x"39a0d315", 
    x"39a0dfb7", 
    x"39a0ec5b", 
    x"39a0f901", 
    x"39a105a9", 
    x"39a11253", 
    x"39a11eff", 
    x"39a12bad", 
    x"39a1385d", 
    x"39a1450f", 
    x"39a151c3", 
    x"39a15e79", 
    x"39a16b31", 
    x"39a177eb", 
    x"39a184a7", 
    x"39a19165", 
    x"39a19e25", 
    x"39a1aae7", 
    x"39a1b7ab", 
    x"39a1c471", 
    x"39a1d13a", 
    x"39a1de04", 
    x"39a1ead0", 
    x"39a1f79e", 
    x"39a2046e", 
    x"39a21140", 
    x"39a21e15", 
    x"39a22aeb", 
    x"39a237c3", 
    x"39a2449e", 
    x"39a2517a", 
    x"39a25e58", 
    x"39a26b39", 
    x"39a2781b", 
    x"39a28500", 
    x"39a291e6", 
    x"39a29ecf", 
    x"39a2abba", 
    x"39a2b8a7", 
    x"39a2c595", 
    x"39a2d286", 
    x"39a2df79", 
    x"39a2ec6e", 
    x"39a2f965", 
    x"39a3065e", 
    x"39a31359", 
    x"39a32057", 
    x"39a32d56", 
    x"39a33a57", 
    x"39a3475b", 
    x"39a35460", 
    x"39a36168", 
    x"39a36e72", 
    x"39a37b7d", 
    x"39a3888b", 
    x"39a3959b", 
    x"39a3a2ad", 
    x"39a3afc1", 
    x"39a3bcd8", 
    x"39a3c9f0", 
    x"39a3d70a", 
    x"39a3e427", 
    x"39a3f145", 
    x"39a3fe66", 
    x"39a40b89", 
    x"39a418ae", 
    x"39a425d5", 
    x"39a432fe", 
    x"39a44029", 
    x"39a44d56", 
    x"39a45a86", 
    x"39a467b7", 
    x"39a474eb", 
    x"39a48221", 
    x"39a48f59", 
    x"39a49c93", 
    x"39a4a9cf", 
    x"39a4b70d", 
    x"39a4c44e", 
    x"39a4d190", 
    x"39a4ded5", 
    x"39a4ec1c", 
    x"39a4f965", 
    x"39a506b0", 
    x"39a513fd", 
    x"39a5214d", 
    x"39a52e9e", 
    x"39a53bf2", 
    x"39a54948", 
    x"39a556a0", 
    x"39a563fa", 
    x"39a57157", 
    x"39a57eb5", 
    x"39a58c16", 
    x"39a59978", 
    x"39a5a6dd", 
    x"39a5b445", 
    x"39a5c1ae", 
    x"39a5cf19", 
    x"39a5dc87", 
    x"39a5e9f7", 
    x"39a5f769", 
    x"39a604dd", 
    x"39a61254", 
    x"39a61fcc", 
    x"39a62d47", 
    x"39a63ac4", 
    x"39a64843", 
    x"39a655c4", 
    x"39a66348", 
    x"39a670cd", 
    x"39a67e55", 
    x"39a68bdf", 
    x"39a6996c", 
    x"39a6a6fa", 
    x"39a6b48b", 
    x"39a6c21e", 
    x"39a6cfb3", 
    x"39a6dd4a", 
    x"39a6eae4", 
    x"39a6f880", 
    x"39a7061e", 
    x"39a713be", 
    x"39a72161", 
    x"39a72f05", 
    x"39a73cac", 
    x"39a74a55", 
    x"39a75801", 
    x"39a765ae", 
    x"39a7735e", 
    x"39a78110", 
    x"39a78ec5", 
    x"39a79c7b", 
    x"39a7aa34", 
    x"39a7b7ef", 
    x"39a7c5ac", 
    x"39a7d36c", 
    x"39a7e12e", 
    x"39a7eef2", 
    x"39a7fcb8", 
    x"39a80a81", 
    x"39a8184c", 
    x"39a82619", 
    x"39a833e8", 
    x"39a841ba", 
    x"39a84f8e", 
    x"39a85d64", 
    x"39a86b3c", 
    x"39a87917", 
    x"39a886f4", 
    x"39a894d3", 
    x"39a8a2b5", 
    x"39a8b099", 
    x"39a8be7f", 
    x"39a8cc68", 
    x"39a8da52", 
    x"39a8e83f", 
    x"39a8f62f", 
    x"39a90420", 
    x"39a91214", 
    x"39a9200b", 
    x"39a92e03", 
    x"39a93bfe", 
    x"39a949fb", 
    x"39a957fb", 
    x"39a965fd", 
    x"39a97401", 
    x"39a98207", 
    x"39a99010", 
    x"39a99e1b", 
    x"39a9ac28", 
    x"39a9ba38", 
    x"39a9c84a", 
    x"39a9d65f", 
    x"39a9e475", 
    x"39a9f28f", 
    x"39aa00aa", 
    x"39aa0ec8", 
    x"39aa1ce8", 
    x"39aa2b0a", 
    x"39aa392f", 
    x"39aa4756", 
    x"39aa5580", 
    x"39aa63ac", 
    x"39aa71da", 
    x"39aa800b", 
    x"39aa8e3e", 
    x"39aa9c73", 
    x"39aaaaab"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
