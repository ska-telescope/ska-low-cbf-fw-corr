-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom2 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom2; 
 
architecture behavioral of inv_rom2 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"3a2ac721", 
    x"3a2ae3a1", 
    x"3a2b002b", 
    x"3a2b1cbe", 
    x"3a2b395a", 
    x"3a2b5601", 
    x"3a2b72b0", 
    x"3a2b8f6a", 
    x"3a2bac2d", 
    x"3a2bc8fa", 
    x"3a2be5d0", 
    x"3a2c02b0", 
    x"3a2c1f9a", 
    x"3a2c3c8d", 
    x"3a2c598b", 
    x"3a2c7692", 
    x"3a2c93a2", 
    x"3a2cb0bd", 
    x"3a2ccde1", 
    x"3a2ceb10", 
    x"3a2d0848", 
    x"3a2d258a", 
    x"3a2d42d6", 
    x"3a2d602b", 
    x"3a2d7d8b", 
    x"3a2d9af5", 
    x"3a2db869", 
    x"3a2dd5e6", 
    x"3a2df36e", 
    x"3a2e1100", 
    x"3a2e2e9b", 
    x"3a2e4c41", 
    x"3a2e69f1", 
    x"3a2e87ab", 
    x"3a2ea570", 
    x"3a2ec33e", 
    x"3a2ee117", 
    x"3a2efefa", 
    x"3a2f1ce7", 
    x"3a2f3ade", 
    x"3a2f58df", 
    x"3a2f76eb", 
    x"3a2f9501", 
    x"3a2fb322", 
    x"3a2fd14c", 
    x"3a2fef82", 
    x"3a300dc1", 
    x"3a302c0b", 
    x"3a304a5f", 
    x"3a3068be", 
    x"3a308727", 
    x"3a30a59b", 
    x"3a30c41a", 
    x"3a30e2a2", 
    x"3a310136", 
    x"3a311fd4", 
    x"3a313e7c", 
    x"3a315d2f", 
    x"3a317bed", 
    x"3a319ab6", 
    x"3a31b989", 
    x"3a31d867", 
    x"3a31f74f", 
    x"3a321643", 
    x"3a323541", 
    x"3a32544a", 
    x"3a32735e", 
    x"3a32927c", 
    x"3a32b1a6", 
    x"3a32d0da", 
    x"3a32f019", 
    x"3a330f63", 
    x"3a332eb8", 
    x"3a334e19", 
    x"3a336d84", 
    x"3a338cfa", 
    x"3a33ac7b", 
    x"3a33cc07", 
    x"3a33eb9e", 
    x"3a340b41", 
    x"3a342aee", 
    x"3a344aa7", 
    x"3a346a6b", 
    x"3a348a3a", 
    x"3a34aa14", 
    x"3a34c9fa", 
    x"3a34e9ea", 
    x"3a3509e7", 
    x"3a3529ee", 
    x"3a354a01", 
    x"3a356a1f", 
    x"3a358a48", 
    x"3a35aa7d", 
    x"3a35cabe", 
    x"3a35eb09", 
    x"3a360b61", 
    x"3a362bc4", 
    x"3a364c32", 
    x"3a366cac", 
    x"3a368d31", 
    x"3a36adc2", 
    x"3a36ce5f", 
    x"3a36ef07", 
    x"3a370fbb", 
    x"3a37307b", 
    x"3a375147", 
    x"3a37721e", 
    x"3a379301", 
    x"3a37b3ef", 
    x"3a37d4ea", 
    x"3a37f5f1", 
    x"3a381703", 
    x"3a383821", 
    x"3a38594b", 
    x"3a387a81", 
    x"3a389bc3", 
    x"3a38bd11", 
    x"3a38de6c", 
    x"3a38ffd2", 
    x"3a392144", 
    x"3a3942c2", 
    x"3a39644d", 
    x"3a3985e3", 
    x"3a39a786", 
    x"3a39c935", 
    x"3a39eaf0", 
    x"3a3a0cb8", 
    x"3a3a2e8c", 
    x"3a3a506c", 
    x"3a3a7258", 
    x"3a3a9451", 
    x"3a3ab656", 
    x"3a3ad868", 
    x"3a3afa86", 
    x"3a3b1cb0", 
    x"3a3b3ee7", 
    x"3a3b612b", 
    x"3a3b837b", 
    x"3a3ba5d7", 
    x"3a3bc841", 
    x"3a3beab6", 
    x"3a3c0d39", 
    x"3a3c2fc8", 
    x"3a3c5264", 
    x"3a3c750d", 
    x"3a3c97c2", 
    x"3a3cba84", 
    x"3a3cdd53", 
    x"3a3d002f", 
    x"3a3d2318", 
    x"3a3d460e", 
    x"3a3d6910", 
    x"3a3d8c20", 
    x"3a3daf3c", 
    x"3a3dd266", 
    x"3a3df59d", 
    x"3a3e18e0", 
    x"3a3e3c31", 
    x"3a3e5f8f", 
    x"3a3e82fa", 
    x"3a3ea672", 
    x"3a3ec9f8", 
    x"3a3eed8b", 
    x"3a3f112b", 
    x"3a3f34d8", 
    x"3a3f5892", 
    x"3a3f7c5b", 
    x"3a3fa030", 
    x"3a3fc413", 
    x"3a3fe803", 
    x"3a400c01", 
    x"3a40300c", 
    x"3a405425", 
    x"3a40784b", 
    x"3a409c7f", 
    x"3a40c0c1", 
    x"3a40e510", 
    x"3a41096d", 
    x"3a412dd8", 
    x"3a415250", 
    x"3a4176d6", 
    x"3a419b6a", 
    x"3a41c00c", 
    x"3a41e4bc", 
    x"3a420979", 
    x"3a422e45", 
    x"3a42531f", 
    x"3a427806", 
    x"3a429cfc", 
    x"3a42c1ff", 
    x"3a42e711", 
    x"3a430c31", 
    x"3a43315f", 
    x"3a43569b", 
    x"3a437be5", 
    x"3a43a13e", 
    x"3a43c6a5", 
    x"3a43ec1a", 
    x"3a44119e", 
    x"3a443730", 
    x"3a445cd0", 
    x"3a44827f", 
    x"3a44a83c", 
    x"3a44ce08", 
    x"3a44f3e2", 
    x"3a4519cb", 
    x"3a453fc2", 
    x"3a4565c8", 
    x"3a458bdd", 
    x"3a45b201", 
    x"3a45d833", 
    x"3a45fe74", 
    x"3a4624c4", 
    x"3a464b22", 
    x"3a467190", 
    x"3a46980c", 
    x"3a46be98", 
    x"3a46e532", 
    x"3a470bdb", 
    x"3a473294", 
    x"3a47595b", 
    x"3a478032", 
    x"3a47a718", 
    x"3a47ce0c", 
    x"3a47f511", 
    x"3a481c24", 
    x"3a484347", 
    x"3a486a79", 
    x"3a4891ba", 
    x"3a48b90b", 
    x"3a48e06b", 
    x"3a4907da", 
    x"3a492f59", 
    x"3a4956e8", 
    x"3a497e86", 
    x"3a49a634", 
    x"3a49cdf1", 
    x"3a49f5bf", 
    x"3a4a1d9b", 
    x"3a4a4588", 
    x"3a4a6d84", 
    x"3a4a9590", 
    x"3a4abdac", 
    x"3a4ae5d8", 
    x"3a4b0e14", 
    x"3a4b3660", 
    x"3a4b5ebc", 
    x"3a4b8728", 
    x"3a4bafa4", 
    x"3a4bd830", 
    x"3a4c00cc", 
    x"3a4c2978", 
    x"3a4c5235", 
    x"3a4c7b02", 
    x"3a4ca3df", 
    x"3a4ccccd", 
    x"3a4cf5cb", 
    x"3a4d1ed9", 
    x"3a4d47f8", 
    x"3a4d7127", 
    x"3a4d9a67", 
    x"3a4dc3b8", 
    x"3a4ded19", 
    x"3a4e168a", 
    x"3a4e400d", 
    x"3a4e69a0", 
    x"3a4e9344", 
    x"3a4ebcf9", 
    x"3a4ee6be", 
    x"3a4f1095", 
    x"3a4f3a7c", 
    x"3a4f6475", 
    x"3a4f8e7e", 
    x"3a4fb899", 
    x"3a4fe2c4", 
    x"3a500d01", 
    x"3a50374f", 
    x"3a5061ae", 
    x"3a508c1e", 
    x"3a50b6a0", 
    x"3a50e133", 
    x"3a510bd7", 
    x"3a51368d", 
    x"3a516154", 
    x"3a518c2d", 
    x"3a51b717", 
    x"3a51e213", 
    x"3a520d21", 
    x"3a523840", 
    x"3a526371", 
    x"3a528eb4", 
    x"3a52ba08", 
    x"3a52e56f", 
    x"3a5310e7", 
    x"3a533c71", 
    x"3a53680d", 
    x"3a5393bb", 
    x"3a53bf7c", 
    x"3a53eb4e", 
    x"3a541733", 
    x"3a544329", 
    x"3a546f32", 
    x"3a549b4d", 
    x"3a54c77b", 
    x"3a54f3bb", 
    x"3a55200d", 
    x"3a554c72", 
    x"3a5578e9", 
    x"3a55a573", 
    x"3a55d210", 
    x"3a55febf", 
    x"3a562b81", 
    x"3a565855", 
    x"3a56853d", 
    x"3a56b237", 
    x"3a56df44", 
    x"3a570c64", 
    x"3a573997", 
    x"3a5766dd", 
    x"3a579436", 
    x"3a57c1a2", 
    x"3a57ef21", 
    x"3a581cb4", 
    x"3a584a5a", 
    x"3a587813", 
    x"3a58a5df", 
    x"3a58d3bf", 
    x"3a5901b2", 
    x"3a592fb9", 
    x"3a595dd3", 
    x"3a598c01", 
    x"3a59ba42", 
    x"3a59e898", 
    x"3a5a1700", 
    x"3a5a457d", 
    x"3a5a740e", 
    x"3a5aa2b2", 
    x"3a5ad16a", 
    x"3a5b0037", 
    x"3a5b2f17", 
    x"3a5b5e0c", 
    x"3a5b8d14", 
    x"3a5bbc31", 
    x"3a5beb62", 
    x"3a5c1aa7", 
    x"3a5c4a01", 
    x"3a5c796f", 
    x"3a5ca8f1", 
    x"3a5cd888", 
    x"3a5d0834", 
    x"3a5d37f4", 
    x"3a5d67c9", 
    x"3a5d97b2", 
    x"3a5dc7b0", 
    x"3a5df7c3", 
    x"3a5e27eb", 
    x"3a5e5828", 
    x"3a5e887a", 
    x"3a5eb8e0", 
    x"3a5ee95c", 
    x"3a5f19ed", 
    x"3a5f4a93", 
    x"3a5f7b4f", 
    x"3a5fac1f", 
    x"3a5fdd05", 
    x"3a600e01", 
    x"3a603f12", 
    x"3a607038", 
    x"3a60a174", 
    x"3a60d2c6", 
    x"3a61042d", 
    x"3a6135aa", 
    x"3a61673d", 
    x"3a6198e5", 
    x"3a61caa4", 
    x"3a61fc78", 
    x"3a622e63", 
    x"3a626063", 
    x"3a62927a", 
    x"3a62c4a7", 
    x"3a62f6ea", 
    x"3a632943", 
    x"3a635bb3", 
    x"3a638e39", 
    x"3a63c0d6", 
    x"3a63f389", 
    x"3a642652", 
    x"3a645933", 
    x"3a648c2a", 
    x"3a64bf38", 
    x"3a64f25d", 
    x"3a652598", 
    x"3a6558eb", 
    x"3a658c54", 
    x"3a65bfd5", 
    x"3a65f36d", 
    x"3a66271c", 
    x"3a665ae2", 
    x"3a668ebf", 
    x"3a66c2b4", 
    x"3a66f6c1", 
    x"3a672ae4", 
    x"3a675f20", 
    x"3a679373", 
    x"3a67c7de", 
    x"3a67fc60", 
    x"3a6830fa", 
    x"3a6865ac", 
    x"3a689a77", 
    x"3a68cf59", 
    x"3a690453", 
    x"3a693965", 
    x"3a696e90", 
    x"3a69a3d2", 
    x"3a69d92d", 
    x"3a6a0ea1", 
    x"3a6a442d", 
    x"3a6a79d1", 
    x"3a6aaf8e", 
    x"3a6ae564", 
    x"3a6b1b52", 
    x"3a6b515a", 
    x"3a6b877a", 
    x"3a6bbdb3", 
    x"3a6bf405", 
    x"3a6c2a70", 
    x"3a6c60f4", 
    x"3a6c9791", 
    x"3a6cce48", 
    x"3a6d0518", 
    x"3a6d3c01", 
    x"3a6d7304", 
    x"3a6daa20", 
    x"3a6de156", 
    x"3a6e18a6", 
    x"3a6e500f", 
    x"3a6e8792", 
    x"3a6ebf2f", 
    x"3a6ef6e6", 
    x"3a6f2eb7", 
    x"3a6f66a2", 
    x"3a6f9ea8", 
    x"3a6fd6c7", 
    x"3a700f01", 
    x"3a704755", 
    x"3a707fc4", 
    x"3a70b84d", 
    x"3a70f0f1", 
    x"3a7129af", 
    x"3a716289", 
    x"3a719b7d", 
    x"3a71d48c", 
    x"3a720db6", 
    x"3a7246fb", 
    x"3a72805b", 
    x"3a72b9d6", 
    x"3a72f36d", 
    x"3a732d1f", 
    x"3a7366ec", 
    x"3a73a0d5", 
    x"3a73dada", 
    x"3a7414fa", 
    x"3a744f36", 
    x"3a74898d", 
    x"3a74c401", 
    x"3a74fe91", 
    x"3a75393c", 
    x"3a757404", 
    x"3a75aee8", 
    x"3a75e9e8", 
    x"3a762505", 
    x"3a76603e", 
    x"3a769b93", 
    x"3a76d705", 
    x"3a771294", 
    x"3a774e40", 
    x"3a778a08", 
    x"3a77c5ee", 
    x"3a7801f0", 
    x"3a783e10", 
    x"3a787a4c", 
    x"3a78b6a6", 
    x"3a78f31d", 
    x"3a792fb2", 
    x"3a796c64", 
    x"3a79a934", 
    x"3a79e622", 
    x"3a7a232d", 
    x"3a7a6056", 
    x"3a7a9d9d", 
    x"3a7adb02", 
    x"3a7b1885", 
    x"3a7b5627", 
    x"3a7b93e6", 
    x"3a7bd1c4", 
    x"3a7c0fc1", 
    x"3a7c4ddc", 
    x"3a7c8c16", 
    x"3a7cca6e", 
    x"3a7d08e5", 
    x"3a7d477b", 
    x"3a7d8631", 
    x"3a7dc505", 
    x"3a7e03f8", 
    x"3a7e430b", 
    x"3a7e823d", 
    x"3a7ec18e", 
    x"3a7f00ff", 
    x"3a7f4090", 
    x"3a7f8040", 
    x"3a7fc010", 
    x"3a800000"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
