----------------------------------------------------------------------------------
-- Company: CSIRO CASS 
-- Engineer: David Humphrey
-- 
-- Create Date: 14.11.2018 11:27:29
-- Module Name: correlatorFBTop25 - Behavioral
-- Description: 
--  Filterbank with 12 FIR taps, 4096 point FFT, critically sampled.
--  Processes 4 parallel signals, each with 8 bit complex data (8 bit real + 8 bit imaginary).
--  This version (with the "25" suffix) refers to the use of 25 bits of precision in the FFT
--  high precision is used to ensure very low bias in the filterbank output (needed to meet the low.CBF 1000 hour noise test).
--  
-- Supporting Code:
--  The Matlab model should be in the directory ../matlab_model
--  Key files:
--   * ../matlab_model/run_correlatorFB.m 
--       Generate input files for the simulation, run the matlab model and compares with simulation output
--   * ../matlab_model/get_rom_coefficients.m
--       Generates ROM data used in the firmware. ROMs are initialised using .coe files.
--       "filtertaps_X.coe" : X runs from 1 to 12, contents of the 12 ROMS used to store the FIR filter taps.
--
--  There is a top level module that can be used to build this in a standalone version 
--   "correlatorFBtesttop.vhd"
-- Structure:
--
--  File Structure
--  --------------
--  Outline of the structure shown below. Excludes .xci files for DSPs, RAMs and ROMs.
--
--    correlatorFBTop.vhd : This file, 4 complex inputs, 12 FIR filter taps, 4096 point FFT.
--        |
--        +-- correlatorFBMem.vhd         : Input memory for the filterbank, 12 blocks of memory chained together. Also holds memory for the coefficients.
--        +-- fb_DSP25.vhd                : 12 TAP FIR filter
--        +-- correlatorFFT25wrapper.vhd  : 4096 point FFT
--                |
--                +-- fft4096_25bit.xci : standard Xilinx 4096 point FFT (4 used).
--
--  TestBench
--  ---------
--  correlatorFB_tb.vhd reads the input data generated by the Matlab model and generates output files for checking by the matlab code.
--
--  Resource Use
--  ------------
--  Approximate resource usage is 
--   LUTs        = 15,607
--   DSPs        = 176
--   Registers   = 27,187
--   BRAMs (36K) = 58
--   URAMs       = 15
--  Note this is about 50% more LUTS and registers as compared with the version that uses 16 bit precision for the FFT (but the same number of DSPs).
-- 
--  Power estimate (Guess based on related measurement on zcu111 board)
--   about 1 W static, 3.5 W dynamic.
--
--  -----------------------------------------------------------------------------------------------
--  Description
--  -----------
--
-- 1. Filterbank Memory
--   The filterbank memory consists of 11 blocks of memory chained together.
--   The read and write addresses are staggered by one clock for each memory, implemented as a 12 sample delay line on
--   the address. This makes the timing easy to meet for the  memory address signals (which would otherwise be high-fanout signals)
--   and also enables use of the adders in the DSPs for the FIR filter.  
--
-- 2. FIR filter
--   The FIR filter uses 12 DSPs for each of the 8 simultaneous samples (4 channels * 2 [real+imaginary]) that are read from the memory.
--   So the FIR filter uses (12 DSPS) * (8 simultaneous samples) = 96 DSPs.
--   The filter is implemented entirely in DSPs. The PCOUT port on the DSP is used to send the result of the multiplication
--   to the next DSP in the chain, where it is added using the adder in the DSP. This scheme requires that the inputs to the
--   12 DSPs are staggered to account for the pipeline stage on the PCOUT port. The staggering is done by controlling the address
--   to the memories as described above.
--
-- 3. 4096 point FFT
--   Standard Xilinx FFT. Some messy logic at the front to account for the delay inserted by the "real-time" mode.
--
-- 4. Reorder memory
--   Data out of the FFT is in bit reversed order. It is stored in a double buffer in order from low to high frequencies,
--   then read out as 3456 fine channels.
----------------------------------------------------------------------------------
library IEEE, common_lib, filterbanks_lib;
use common_lib.common_pkg.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity correlatorFBTop25 is
    generic(
        METABITS : integer := 64;     -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP : integer := 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    );
    port(
        -- clock, target is 380 MHz
        clk : in std_logic;
        rst : in std_logic;
        -- Data input, common valid signal, expects packets of 4096 samples. Requires at least 2 clocks idle time between packets.
        data0_i : in t_slv_16_arr(1 downto 0);  -- 4 Inputs, each complex data, 16 bit real, 16 bit imaginary.
        data1_i : in t_slv_16_arr(1 downto 0);
        data2_i : in t_slv_16_arr(1 downto 0);
        data3_i : in t_slv_16_arr(1 downto 0);
        RFI_threshold01_i : in std_logic_vector(31 downto 0);
        RFI_threshold23_i : in std_logic_vector(31 downto 0);
        meta_i  : in std_logic_vector((METABITS-1) downto 0);
        valid_i : in std_logic;
        -- Data out; bursts of 3456 clocks for each channel.
        data0_o : out t_slv_16_arr(1 downto 0);   -- 4 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o : out t_slv_16_arr(1 downto 0);
        data2_o : out t_slv_16_arr(1 downto 0);
        data3_o : out t_slv_16_arr(1 downto 0);
        meta_o  : out std_logic_vector((METABITS-1) downto 0);
        mark_RFI01_o : out std_logic;
        mark_RFI23_o : out std_logic;
        valid_o : out std_logic;
        -- Writing FIR Taps
        FIRTapData_i : in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i : in std_logic_vector(15 downto 0);  -- 4096 * 12 filter taps = 49152 total.
        FIRTapWE_i   : in std_logic;
        FIRTapClk    : in std_logic
    );
end correlatorFBTop25;

architecture Behavioral of correlatorFBTop25 is
    
    signal wrData128 : std_logic_vector(127 downto 0);
    signal FBmemRdData : t_slv_128_arr(11 downto 0);
    signal FBmemFIRTaps, FBmemFIRTapsDel : t_slv_18_arr(11 downto 0);
    
    type fbtype is array(7 downto 0) of t_slv_16_arr(11 downto 0);
    signal FBRdData, FBRdDataDel : fbtype; 
    signal FIRDout : t_slv_25_arr(7 downto 0);
    signal fftIndex : t_slv_12_arr(3 downto 0);
    
    signal fftRealOut : t_slv_16_arr(3 downto 0);
    signal fftImagOut : t_slv_16_arr(3 downto 0);
    signal fftvalidOut : std_logic_vector(3 downto 0) := "0000";
    
    signal startAdv : std_logic_vector(31 downto 0);
    signal validDel1, validDel2, validDel3 : std_logic := '0';
    signal startFFT : std_logic := '0';
    
    signal reorderDout0, reorderDout1, reorderDout2, reorderDout3 : std_logic_vector(63 downto 0);
    signal reorderWE : std_logic_vector(1 downto 0);
    signal reorderWrAddr : std_logic_vector(11 downto 0);
    signal reorderRdAddr : std_logic_vector(11 downto 0);
    signal bufSelectWr, bufSelectRd : std_logic := '0';
    signal reorderDin0, reorderDin1 : std_logic_vector(63 downto 0);
    signal rdRunning : std_logic := '0';
    signal rdRunningDel2, rdRunningDel1 : std_logic := '0';
    signal validOutDel1 : std_logic := '0';
    signal bufSelectRdDel1, bufSelectRdDel2 : std_logic := '0';
    
    signal metaDel0, metaDel1, metaDel2, metaDel3, metaDel4 : std_logic_vector(METABITS+16-1 downto 0);
    signal metaOut : std_logic_vector((METABITS-1) downto 0);
    signal outputCountOut : std_logic_vector(15 downto 0);
    signal outputCount : std_logic_vector(15 downto 0);
    signal metaDel1Count, metaDel2Count, metaDel3Count : std_logic_vector(11 downto 0);
    signal FBmemRdAddr : t_slv_12_arr(11 downto 0);
    
    signal RFI_flagged : t_slv_12_arr(1 downto 0);
    signal RFI_count_start, RFI_count_last, RFI_count_last_del1 : std_logic_vector(11 downto 0) := "000000000000";
    type RFI_sum_type is array(1 downto 0) of t_slv_10_arr(11 downto 0);
    signal RFI_sum, RFI_sum_store : RFI_sum_type;
    signal RFI_count_1024block_del1, RFI_count_1024block : std_logic_vector(2 downto 0);
    signal RFI_weight_addr, RFI_weight_addr_del1, RFI_weight_addr_del2 : std_logic_vector(6 downto 0);
    signal RFI_weight_addr_low : std_logic_vector(2 downto 0);
    signal RFI_weight_FIR_tap : std_logic_vector(3 downto 0);
    signal mark_as_RFI23_del2, mark_as_RFI23_del1, mark_as_RFI01_del2, mark_as_RFI01_del1 : std_logic := '0';
    type RFI_fsm_type is  (run, check_threshold, idle);
    signal RFI_fsm, RFI_fsm_del1, RFI_fsm_del2 : RFI_fsm_type := idle;
    signal RFI_sum_station0, RFI_sum_station1 : std_logic_vector(9 downto 0);
    signal RFI_sum_station0_ext, RFI_sum_station1_ext : std_logic_vector(10 downto 0);
    signal RFI_weighted_sum0, RFI_weighted_sum1 : signed(32 downto 0);
    signal RFI_weighted_sum0_ext, RFI_weighted_sum1_ext : std_logic_vector(39 downto 0);
    signal final_RFI_sum0, final_RFI_sum1 : std_logic_vector(39 downto 0);
    signal mark_as_RFI01, mark_as_RFI23 : std_logic := '0';
    signal mark_as_RFI_valid : std_logic := '0';
    signal RFI_weight : std_logic_vector(21 downto 0);
    signal RFI_threshold01_max, RFI_threshold23_max : std_logic := '0';
    signal RFI_threshold01_hold, RFI_threshold23_hold, RFI_threshold23_del1, RFI_threshold01_del1 : std_logic_vector(31 downto 0) := (others => '0');
    
begin
    
    ------------------------------------------------------------------------------------
    -- 1. Input Memory
    -- ---------------
    
    wrData128 <= data3_i(1) & data3_i(0) & data2_i(1) & data2_i(0) & data1_i(1) & data1_i(0) & data0_i(1) & data0_i(0);

    cmem : entity filterbanks_lib.correlatorFBMem
    generic map (
        TAPS => 12)  -- Note only partially parameterized; modification needed to support anything other than 12.
    port map (
        clk      => clk,
        -- Write data for the start of the chain
        wrData_i => wrData128,        -- in(127:0);
        wrEn_i   => valid_i,          -- in std_logic; should be a burst of 4096 clocks.
        -- Read data, comes out 2 clocks after the first write.
        rd_data_o  => FBmemRdData,    -- out t_slv_128_arr(TAPS-1 downto 0); 64 bits wide, 12 taps simultaneously; First sample is wr_data_i delayed by 1 clock. 
        rd_data_addr_o => FBmemRdAddr, -- out t_slv_12_arr(TAPS-1 downto 0); The address (0 to 4095) that the corresponding data in rd_data_o comes from
        coef_o     => FBmemFIRTaps,   -- out t_slv_18_arr(TAPS-1 downto 0);  18 bits per filter tap.
        -- Writing FIR Taps
        FIRTapData_i => FIRTapData_i, -- in(17:0);  -- For register writes of the filtertaps.
        FIRTapData_o => FIRTapData_o, -- out(17:0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i => FIRTapAddr_i, -- in(15:0);  -- 4096 * 12 filter taps = 49152 total.
        FIRTapWE_i   => FIRTapWE_i,   -- in std_logic;
        FIRTapClk    => FIRTapClk     -- in std_logic
    );


    -------------------------------------------------------------------------------------
    -- 2. FIR filter
    -- -------------
    -- 8 instances, 4 channels * (real + imaginary). Same filter taps used for all.
    -- In low.CBF, processes simultaneously 2 (real+imaginary) * 2 (stations) * 2 (polarisations) = 8
    -- 
    
    CsampleGen : for j in 0 to 7 generate
        coefGen : for k in 0 to 11 generate
            FBRdData(j)(k) <= FBmemRdData(k)((j*16 + 15) downto (j*16));
        end generate;
    end generate;
    
    -- Extra pipeline stage so that BRAMs and URAMs can be placed further from the DSP.
    -- (without this pipeline stage, the output register in the URAM connects to the input register in the DSP).
    -- Also calculate the RFI metrics
    process(clk)
    begin
        if rising_edge(clk) then
            FBmemFIRTapsDel <= FBmemFIRTaps;
            
            -- Accumulate the number of RFI flagged samples in each 512 sample block
            for j in 0 to 1 loop
                -- j indexes the station; 4 streams per station (2 pol x (re+im)), if any of the 4 samples are flagged then all are flagged.
                for k in 0 to 11 loop
                    -- pipeline stage to identify flagged samples
                    if FBRdData(j*4 + 0)(k) = x"8000" or FBRdData(j*4 + 1)(k) = x"8000" or FBRdData(j*4 + 2)(k) = x"8000" or FBRdData(j*4 + 3)(k) = x"8000" then
                        RFI_flagged(j)(k) <= '1';
                    else
                        RFI_flagged(j)(k) <= '0';
                    end if;
                    -- Accumulate the number of flagged samples across every 512 samples
                    if RFI_count_start(k) = '1' then
                        -- This is the first sample in a block of 512 samples
                        if RFI_flagged(j)(k) = '1' then
                            RFI_sum(j)(k) <= "0000000001";
                        else
                            RFI_sum(j)(k) <= "0000000000";
                        end if;
                    elsif RFI_flagged(j)(k) = '1' then
                        RFI_sum(j)(k) <= std_logic_vector(unsigned(RFI_sum(j)(k)) + 1);
                    end if;
                    -- Store RFI counts for processing
                    if RFI_count_last_del1(k) = '1' then
                        RFI_sum_store(j)(k) <= RFI_sum(j)(k);
                    end if;
                end loop;
            end loop;

            for k in 0 to 11 loop
                if FBmemRdAddr(k)(8 downto 0) = "000000000" then
                    -- Start of every 512 sample block
                    RFI_count_start(k) <= '1';
                else
                    RFI_count_start(k) <= '0';
                end if;
                if FBmemRdAddr(k)(8 downto 0) = "111111111" then 
                    RFI_count_last(k) <= '1';
                else
                    RFI_count_last(k) <= '0';
                end if;
            end loop;
            RFI_count_last_del1 <= RFI_count_last;        

            if FBmemRdAddr(11)(8 downto 0) = "111111111" then
                RFI_count_1024block <= FBmemRdAddr(11)(11 downto 9);
            end if;
            RFI_count_1024block_del1 <= RFI_count_1024block;
            
            -- 
            if RFI_count_last_del1(11) = '1' then
                RFI_fsm <= run;
                RFI_weight_addr_low <= RFI_count_1024block_del1;
                RFI_weight_FIR_tap <= "0000";
            else
                case RFI_fsm is
                    when run =>
                        -- Go through all 12 counts in RFI_sum_store, weight them and sum 
                        -- to get an estimate of the total error in the output 
                        if unsigned(RFI_weight_FIR_tap) = 11 then
                            if RFI_weight_addr_low = "111" then
                                -- final sum complete, compare with the allowed threshold
                                RFI_fsm <= check_threshold;
                            else
                                RFI_fsm <= idle;
                            end if;
                        end if;
                        RFI_weight_FIR_tap <= std_logic_vector(unsigned(RFI_weight_FIR_tap) + 1);
                    
                    when check_threshold =>
                        RFI_fsm <= idle;
                    
                    when idle =>
                        RFI_fsm <= idle;
                    
                    when others =>
                        RFI_fsm <= idle;
                end case;
            end if;
            
            -- case statement since it only runs to 11, and simulation falls over when 
            -- the index (RFI_weight_FIR_tap) is 12.
            case RFI_weight_FIR_tap is
                when "0000" => 
                    RFI_sum_station0 <= RFI_sum_store(0)(0); -- 10 bit value, maximum possible is 512
                    RFI_sum_station1 <= RFI_sum_store(1)(0);
                when "0001" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(1);
                    RFI_sum_station1 <= RFI_sum_store(1)(1);
                when "0010" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(2);
                    RFI_sum_station1 <= RFI_sum_store(1)(2);
                when "0011" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(3);
                    RFI_sum_station1 <= RFI_sum_store(1)(3);
                when "0100" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(4);
                    RFI_sum_station1 <= RFI_sum_store(1)(4);
                when "0101" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(5);
                    RFI_sum_station1 <= RFI_sum_store(1)(5);
                when "0110" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(6);
                    RFI_sum_station1 <= RFI_sum_store(1)(6);
                when "0111" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(7);
                    RFI_sum_station1 <= RFI_sum_store(1)(7);
                when "1000" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(8);
                    RFI_sum_station1 <= RFI_sum_store(1)(8);
                when "1001" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(9);
                    RFI_sum_station1 <= RFI_sum_store(1)(9);
                when "1010" =>
                    RFI_sum_station0 <= RFI_sum_store(0)(10);
                    RFI_sum_station1 <= RFI_sum_store(1)(10);
                when others =>
                    RFI_sum_station0 <= RFI_sum_store(0)(11);
                    RFI_sum_station1 <= RFI_sum_store(1)(11);
            end case;
                
            RFI_weight_addr_del1 <= RFI_weight_addr;
            RFI_fsm_del1 <= RFI_fsm;
            
            RFI_weighted_sum0 <= signed(RFI_sum_station0_ext) * signed(RFI_weight); -- 11 bit x 22 bit = 33 bit result
            RFI_weighted_sum1 <= signed(RFI_sum_station1_ext) * signed(RFI_weight);
            RFI_weight_addr_del2 <= RFI_weight_addr_del1;
            RFI_fsm_del2 <= RFI_fsm_del1;
            
            if RFI_weight_addr_del2 = "0000000" and (RFI_fsm_del2 = run) then
                -- First RFI sum to accumulate
                final_RFI_sum0 <= "0000000" & std_logic_vector(RFI_weighted_sum0);
                final_RFI_sum1 <= "0000000" & std_logic_vector(RFI_weighted_sum1);
            elsif RFI_fsm_del2 = run then
                -- Accumulate
                final_RFI_sum0 <= std_logic_vector(unsigned(final_RFI_sum0) + unsigned(RFI_weighted_sum0_ext));
                final_RFI_sum1 <= std_logic_vector(unsigned(final_RFI_sum1) + unsigned(RFI_weighted_sum1_ext));
            end if;
            
            RFI_threshold01_del1 <= RFI_threshold01_i;
            RFI_threshold23_del1 <= RFI_threshold23_i;
            if valid_i = '0' and validDel1 = '1' then 
                -- On the falling edge of valid, hold the RFI threshold for use a short time later 
                RFI_threshold01_hold <= RFI_threshold01_del1;
                RFI_threshold23_hold <= RFI_threshold23_del1;
            end if;
            
            if RFI_threshold01_hold = x"ffffffff" then 
                RFI_threshold01_max <= '1';
            else
                RFI_threshold01_max <= '0';
            end if;
            
            if RFI_threshold23_hold = x"ffffffff" then 
                RFI_threshold23_max <= '1';
            else
                RFI_threshold23_max <= '0';
            end if;
            
            if RFI_fsm_del2 = check_threshold then
                if ((unsigned(final_RFI_sum0) > unsigned(RFI_threshold01_hold)) and RFI_threshold01_max = '0') then
                    mark_as_RFI01 <= '1';
                else
                    mark_as_RFI01 <= '0';
                end if;
                if ((unsigned(final_RFI_sum1) > unsigned(RFI_threshold23_hold)) and RFI_threshold23_max = '0') then
                    mark_as_RFI23 <= '1';
                else
                    mark_as_RFI23 <= '0';
                end if;
                mark_as_RFI_valid <= '1';
            else
                mark_as_RFI_valid <= '0';
            end if;
            
            -- Replace RFI marked samples with zeros for processing through the filterbank
            for j in 0 to 7 loop
                for k in 0 to 11 loop
                    if FBRdData(j)(k) = x"8000" then
                        FBRdDataDel(j)(k) <= x"0000";
                    else
                        FBRdDataDel(j)(k) <= FBRdData(j)(k);
                    end if;
                end loop;
            end loop;
            
        end if;
    end process;
    
    RFI_sum_station0_ext <= '0' & RFI_sum_station0; -- sign extend so it can be treated as a signed value in the multiply
    RFI_sum_station1_ext <= '0' & RFI_sum_station1;
    
    RFI_weighted_sum0_ext <= "0000000" & std_logic_vector(RFI_weighted_sum0);
    RFI_weighted_sum1_ext <= "0000000" & std_logic_vector(RFI_weighted_sum1);
    
    RFI_weight_addr(2 downto 0) <= RFI_weight_addr_low;
    RFI_weight_addr(6 downto 3) <= RFI_weight_FIR_tap;
    
    RFI_weights_romi : entity filterbanks_lib.RFI_weights
    port map (
        clk    => clk,
        -- 6 bit address
        -- low 2 bits selects the block of 1024 within each block of 4096
        -- High 4 bits selects the FIR tap, valid range 0 to 11
        i_addr => RFI_weight_addr, -- in (6:0)
        -- 1 cycle read latency from i_addr
        o_RFI_weight => RFI_weight  -- out (21:0); 22 bit average RFI-induced power for samples in this block of 512 FIR samples
    );
    
    sampleGen : for j in 0 to 7 generate
            
        FIR : entity filterbanks_lib.fb_DSP25
        generic map (
            TAPS => 12)  -- The module instantiates this number of DSPs
        port map (
            clk    => clk,
            data_i => FBRdDataDel(j),  -- in t_slv_16_arr(11 downto 0);
            coef_i => FBmemFIRTapsDel, -- in t_slv_18_arr(11 downto 0);
            data_o => FIRDout(j)    -- out(24:0)
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 3. FFT
    -- -----------------
    -- 4 x 4096 point FFTs.
    
    process(clk)
    begin
        if rising_edge(clk) then
            validDel1 <= valid_i;
            validDel2 <= validDel1;
            validDel3 <= validDel2;
            if validDel2 = '1' and validDel3 = '0' then
                startAdv(0) <= '1';
            else
                startAdv(0) <= '0';
            end if;
            
            startAdv(31 downto 1) <= startAdv(30 downto 0);
            startFFT <= startAdv(12); -- Delay accounts for the delay through the FIR filter 
            
            -- meta and output count
            -- Once a packet comes it data comes out after a fixed latency, but the gap between packets is variable.
            -- So we use a delay line which shifts after 4095 clocks if there is data in it. 
            if rst = '1' then
                outputCount <= (others => '0'); -- count of the number of packets, used to drop the first 11 output packets.
            elsif valid_i = '1' and validDel1 = '0' then -- rising edge of valid
                outputCount <= std_logic_vector(unsigned(outputCount) + 1);
                metaDel0 <= outputCount & meta_i;
            end if;
            
            if valid_i = '0' and validDel1 = '1' then -- falling edge of valid
                metaDel1 <= metaDel0;
                metaDel1Count <= "111111111111";
            elsif metaDel1Count /= "000000000000" then
                metaDel1Count <= std_logic_vector(unsigned(metaDel1Count) - 1);
            end if;
            
            if mark_as_RFI_valid = '1' then -- occurs about 8 clocks after falling edge of valid_i
                mark_as_RFI01_del1 <= mark_as_RFI01;
                mark_as_RFI23_del1 <= mark_as_RFI23;
            end if;
            
            if metaDel1Count = "000000000001" then
                metaDel2 <= metaDel1;
                mark_as_RFI01_del2 <= mark_as_RFI01_del1;
                mark_as_RFI23_del2 <= mark_as_RFI23_del1;
                metaDel2Count <= "111111111111";
            elsif metaDel2Count /= "000000000000" then
                metaDel2Count <= std_logic_vector(unsigned(metaDel2Count) - 1);
            end if;
            
            if metaDel2Count = "000000000001" then
                metaDel3 <= metaDel2;
                metaDel3Count <= "111111111111";
            elsif metaDel3Count /= "000000000000" then
                metaDel3Count <= std_logic_vector(unsigned(metaDel3Count) - 1);
            end if;
            
            if metaDel3Count = "000000000001" then
                metaDel4 <= metaDel3;
            end if;
            
        end if;
    end process;
    
    
    fftgen : for j in 0 to 3 generate
        
        fft4096 : entity filterbanks_lib.correlatorFFT25wrapper
        port map (
            clk  => clk,
            -- Input
            real_i  => FIRDout(j*2),     -- in(24:0); -- 25 bit real data
            imag_i  => FIRDout(j*2 + 1), -- in(24:0); -- 25 bit imaginary data
            start_i => startFFT,         -- in std_logic;                     -- pulse high; one clock in advance of the data ?
            -- Output
            real_o  => fftRealOut(j), -- out(15:0);
            imag_o  => fftImagOut(j), -- out(15:0);
            index_o => fftIndex(j),   -- out(11:0);
            valid_o => fftvalidOut(j) -- out std_logic
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 4. Reorder the output from bit-reversed to the central 3456 channels, low to high frequency. 
    -- 
    -- Uses an ultraRAM double buffer.
      
    process(clk)
    begin
        if rising_edge(clk) then
        
            if (fftvalidOut(0) = '1' and (signed(fftIndex(0)) > -1729) and (signed(fftIndex(0)) < 1728)) then
                if bufSelectWr = '0' then
                    reorderWE(0) <= '1';
                    reorderWE(1) <= '0';
                else
                    reorderWE(0) <= '0';
                    reorderWE(1) <= '1';
                end if;
            else
                reorderWE(0) <= '0';
                reorderWE(1) <= '0';
            end if;
            reorderWrAddr <= std_logic_vector(signed(fftIndex(0)) + 1728);
            reorderDin0 <= fftImagOut(1) & fftRealOut(1) & fftImagOut(0) & fftRealOut(0);
            reorderDin1 <= fftImagOut(3) & fftRealOut(3) & fftImagOut(2) & fftRealOut(2);
            
            -- Falling edge of validOut triggers reading of the data from the memory
            validOutDel1 <= fftvalidOut(0);
            if fftvalidOut(0) = '0' and validOutDel1 = '1' then
                reorderRdAddr <= "000000000000";
                bufSelectWr <= not bufSelectWr;
                bufSelectRd <= bufSelectWr;
                rdRunning <= '1';
            elsif rdRunning = '1' then
                reorderRdAddr <= std_logic_vector(unsigned(reorderRdAddr) + 1);
                -- read address runs from 0 to 3455
                if unsigned(reorderRdAddr) = 3455 then
                   rdRunning <= '0';
                end if;
            end if;
            rdRunningDel1 <= rdRunning;
            rdRunningDel2 <= rdRunningDel1;
            bufSelectRdDel1 <= bufSelectRd;
            bufSelectRdDel2 <= bufSelectRdDel1;
        end if;
    end process;

    -- Two URAMs for first half of the double buffer
    reorderURAM0 : entity filterbanks_lib.URAM64wrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin0,   -- in(63:0);
        we     => reorderWE(0),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout0   -- out(63:0)
    );

    reorderURAM1 : entity filterbanks_lib.URAM64wrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin1,   -- in(63:0);
        we     => reorderWE(0),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout1   -- out(63:0)
    );    
    
    -- Two URAMs for the second half of the double buffer
    reorderURAM2 : entity filterbanks_lib.URAM64wrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin0,   -- in(63:0);
        we     => reorderWE(1),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout2   -- out(63:0)
    );

    reorderURAM3 : entity filterbanks_lib.URAM64wrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin1,   -- in(63:0);
        we     => reorderWE(1),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout3   -- out(63:0)
    );    
    

    process(clk)
    begin
        if rising_edge(clk) then
            if rdRunningDel1 = '1' and rdRunningDel2 = '0' then -- Rising edge of rdRunning, two clocks prior to valid_o
                metaOut <= metaDel2((METABITS-1) downto 0);
                mark_RFI01_o <= mark_as_RFI01_del2;
                mark_RFI23_o <= mark_as_RFI23_del2;
                outputCountOut <= metaDel2((METABITS+15) downto METABITS);
            end if;
            
            if bufSelectRdDel2 = '0' then
                data0_o(0) <= reorderDout0(15 downto 0);
                data0_o(1) <= reorderDout0(31 downto 16);
                data1_o(0) <= reorderDout0(47 downto 32);
                data1_o(1) <= reorderDout0(63 downto 48);
                data2_o(0) <= reorderDout1(15 downto 0);
                data2_o(1) <= reorderDout1(31 downto 16);
                data3_o(0) <= reorderDout1(47 downto 32);
                data3_o(1) <= reorderDout1(63 downto 48);
            else
                data0_o(0) <= reorderDout2(15 downto 0);
                data0_o(1) <= reorderDout2(31 downto 16);
                data1_o(0) <= reorderDout2(47 downto 32);
                data1_o(1) <= reorderDout2(63 downto 48);
                data2_o(0) <= reorderDout3(15 downto 0);
                data2_o(1) <= reorderDout3(31 downto 16);
                data3_o(0) <= reorderDout3(47 downto 32);
                data3_o(1) <= reorderDout3(63 downto 48);
            end if;
            
            -- outputCountOut counts output packets, starting from 0.
            if (unsigned(outputCountOut) >= FRAMESTODROP) then
                valid_o <= rdRunningDel2;
            else
                valid_o <= '0';
            end if;
            
        end if;
    end process;    
    
    meta_o <= metaOut;
    
end Behavioral;
