-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom4 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom4; 
 
architecture behavioral of inv_rom4 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"3a000000", 
    x"39ffe004", 
    x"39ffc010", 
    x"39ffa024", 
    x"39ff8040", 
    x"39ff6064", 
    x"39ff4090", 
    x"39ff20c3", 
    x"39ff00ff", 
    x"39fee143", 
    x"39fec18e", 
    x"39fea1e1", 
    x"39fe823d", 
    x"39fe62a0", 
    x"39fe430b", 
    x"39fe237d", 
    x"39fe03f8", 
    x"39fde47a", 
    x"39fdc505", 
    x"39fda597", 
    x"39fd8631", 
    x"39fd66d2", 
    x"39fd477b", 
    x"39fd282d", 
    x"39fd08e5", 
    x"39fce9a6", 
    x"39fcca6e", 
    x"39fcab3e", 
    x"39fc8c16", 
    x"39fc6cf5", 
    x"39fc4ddc", 
    x"39fc2ecb", 
    x"39fc0fc1", 
    x"39fbf0bf", 
    x"39fbd1c4", 
    x"39fbb2d2", 
    x"39fb93e6", 
    x"39fb7503", 
    x"39fb5627", 
    x"39fb3752", 
    x"39fb1885", 
    x"39faf9c0", 
    x"39fadb02", 
    x"39fabc4c", 
    x"39fa9d9d", 
    x"39fa7ef6", 
    x"39fa6056", 
    x"39fa41be", 
    x"39fa232d", 
    x"39fa04a4", 
    x"39f9e622", 
    x"39f9c7a7", 
    x"39f9a934", 
    x"39f98ac9", 
    x"39f96c64", 
    x"39f94e08", 
    x"39f92fb2", 
    x"39f91164", 
    x"39f8f31d", 
    x"39f8d4de", 
    x"39f8b6a6", 
    x"39f89876", 
    x"39f87a4c", 
    x"39f85c2a", 
    x"39f83e10", 
    x"39f81ffc", 
    x"39f801f0", 
    x"39f7e3eb", 
    x"39f7c5ee", 
    x"39f7a7f7", 
    x"39f78a08", 
    x"39f76c20", 
    x"39f74e40", 
    x"39f73066", 
    x"39f71294", 
    x"39f6f4c9", 
    x"39f6d705", 
    x"39f6b949", 
    x"39f69b93", 
    x"39f67de5", 
    x"39f6603e", 
    x"39f6429e", 
    x"39f62505", 
    x"39f60773", 
    x"39f5e9e8", 
    x"39f5cc64", 
    x"39f5aee8", 
    x"39f59172", 
    x"39f57404", 
    x"39f5569c", 
    x"39f5393c", 
    x"39f51be3", 
    x"39f4fe91", 
    x"39f4e145", 
    x"39f4c401", 
    x"39f4a6c4", 
    x"39f4898d", 
    x"39f46c5e", 
    x"39f44f36", 
    x"39f43214", 
    x"39f414fa", 
    x"39f3f7e6", 
    x"39f3dada", 
    x"39f3bdd4", 
    x"39f3a0d5", 
    x"39f383dd", 
    x"39f366ec", 
    x"39f34a02", 
    x"39f32d1f", 
    x"39f31042", 
    x"39f2f36d", 
    x"39f2d69e", 
    x"39f2b9d6", 
    x"39f29d15", 
    x"39f2805b", 
    x"39f263a7", 
    x"39f246fb", 
    x"39f22a55", 
    x"39f20db6", 
    x"39f1f11d", 
    x"39f1d48c", 
    x"39f1b801", 
    x"39f19b7d", 
    x"39f17eff", 
    x"39f16289", 
    x"39f14619", 
    x"39f129af", 
    x"39f10d4d", 
    x"39f0f0f1", 
    x"39f0d49c", 
    x"39f0b84d", 
    x"39f09c05", 
    x"39f07fc4", 
    x"39f06389", 
    x"39f04755", 
    x"39f02b28", 
    x"39f00f01", 
    x"39eff2e1", 
    x"39efd6c7", 
    x"39efbab4", 
    x"39ef9ea8", 
    x"39ef82a2", 
    x"39ef66a2", 
    x"39ef4aa9", 
    x"39ef2eb7", 
    x"39ef12cb", 
    x"39eef6e6", 
    x"39eedb07", 
    x"39eebf2f", 
    x"39eea35d", 
    x"39ee8792", 
    x"39ee6bcd", 
    x"39ee500f", 
    x"39ee3457", 
    x"39ee18a6", 
    x"39edfcfb", 
    x"39ede156", 
    x"39edc5b8", 
    x"39edaa20", 
    x"39ed8e8f", 
    x"39ed7304", 
    x"39ed577f", 
    x"39ed3c01", 
    x"39ed2089", 
    x"39ed0518", 
    x"39ece9ac", 
    x"39ecce48", 
    x"39ecb2e9", 
    x"39ec9791", 
    x"39ec7c3f", 
    x"39ec60f4", 
    x"39ec45af", 
    x"39ec2a70", 
    x"39ec0f37", 
    x"39ebf405", 
    x"39ebd8d9", 
    x"39ebbdb3", 
    x"39eba293", 
    x"39eb877a", 
    x"39eb6c67", 
    x"39eb515a", 
    x"39eb3653", 
    x"39eb1b52", 
    x"39eb0058", 
    x"39eae564", 
    x"39eaca76", 
    x"39eaaf8e", 
    x"39ea94ad", 
    x"39ea79d1", 
    x"39ea5efc", 
    x"39ea442d", 
    x"39ea2964", 
    x"39ea0ea1", 
    x"39e9f3e4", 
    x"39e9d92d", 
    x"39e9be7d", 
    x"39e9a3d2", 
    x"39e9892e", 
    x"39e96e90", 
    x"39e953f7", 
    x"39e93965", 
    x"39e91ed9", 
    x"39e90453", 
    x"39e8e9d3", 
    x"39e8cf59", 
    x"39e8b4e5", 
    x"39e89a77", 
    x"39e8800f", 
    x"39e865ac", 
    x"39e84b50", 
    x"39e830fa", 
    x"39e816aa", 
    x"39e7fc60", 
    x"39e7e21c", 
    x"39e7c7de", 
    x"39e7ada5", 
    x"39e79373", 
    x"39e77946", 
    x"39e75f20", 
    x"39e744ff", 
    x"39e72ae4", 
    x"39e710d0", 
    x"39e6f6c1", 
    x"39e6dcb8", 
    x"39e6c2b4", 
    x"39e6a8b7", 
    x"39e68ebf", 
    x"39e674ce", 
    x"39e65ae2", 
    x"39e640fc", 
    x"39e6271c", 
    x"39e60d41", 
    x"39e5f36d", 
    x"39e5d99e", 
    x"39e5bfd5", 
    x"39e5a612", 
    x"39e58c54", 
    x"39e5729d", 
    x"39e558eb", 
    x"39e53f3f", 
    x"39e52598", 
    x"39e50bf8", 
    x"39e4f25d", 
    x"39e4d8c7", 
    x"39e4bf38", 
    x"39e4a5ae", 
    x"39e48c2a", 
    x"39e472ac", 
    x"39e45933", 
    x"39e43fc0", 
    x"39e42652", 
    x"39e40ceb", 
    x"39e3f389", 
    x"39e3da2c", 
    x"39e3c0d6", 
    x"39e3a784", 
    x"39e38e39", 
    x"39e374f3", 
    x"39e35bb3", 
    x"39e34278", 
    x"39e32943", 
    x"39e31014", 
    x"39e2f6ea", 
    x"39e2ddc5", 
    x"39e2c4a7", 
    x"39e2ab8d", 
    x"39e2927a", 
    x"39e2796c", 
    x"39e26063", 
    x"39e24760", 
    x"39e22e63", 
    x"39e2156b", 
    x"39e1fc78", 
    x"39e1e38b", 
    x"39e1caa4", 
    x"39e1b1c2", 
    x"39e198e5", 
    x"39e1800e", 
    x"39e1673d", 
    x"39e14e70", 
    x"39e135aa", 
    x"39e11ce9", 
    x"39e1042d", 
    x"39e0eb77", 
    x"39e0d2c6", 
    x"39e0ba1a", 
    x"39e0a174", 
    x"39e088d3", 
    x"39e07038", 
    x"39e057a2", 
    x"39e03f12", 
    x"39e02687", 
    x"39e00e01", 
    x"39dff580", 
    x"39dfdd05", 
    x"39dfc490", 
    x"39dfac1f", 
    x"39df93b4", 
    x"39df7b4f", 
    x"39df62ee", 
    x"39df4a93", 
    x"39df323e", 
    x"39df19ed", 
    x"39df01a2", 
    x"39dee95c", 
    x"39ded11c", 
    x"39deb8e0", 
    x"39dea0aa", 
    x"39de887a", 
    x"39de704e", 
    x"39de5828", 
    x"39de4007", 
    x"39de27eb", 
    x"39de0fd5", 
    x"39ddf7c3", 
    x"39dddfb7", 
    x"39ddc7b0", 
    x"39ddafaf", 
    x"39dd97b2", 
    x"39dd7fbb", 
    x"39dd67c9", 
    x"39dd4fdc", 
    x"39dd37f4", 
    x"39dd2011", 
    x"39dd0834", 
    x"39dcf05b", 
    x"39dcd888", 
    x"39dcc0ba", 
    x"39dca8f1", 
    x"39dc912e", 
    x"39dc796f", 
    x"39dc61b5", 
    x"39dc4a01", 
    x"39dc3251", 
    x"39dc1aa7", 
    x"39dc0302", 
    x"39dbeb62", 
    x"39dbd3c7", 
    x"39dbbc31", 
    x"39dba4a0", 
    x"39db8d14", 
    x"39db758d", 
    x"39db5e0c", 
    x"39db468f", 
    x"39db2f17", 
    x"39db17a4", 
    x"39db0037", 
    x"39dae8ce", 
    x"39dad16a", 
    x"39daba0c", 
    x"39daa2b2", 
    x"39da8b5d", 
    x"39da740e", 
    x"39da5cc3", 
    x"39da457d", 
    x"39da2e3c", 
    x"39da1700", 
    x"39d9ffca", 
    x"39d9e898", 
    x"39d9d16a", 
    x"39d9ba42", 
    x"39d9a31f", 
    x"39d98c01", 
    x"39d974e7", 
    x"39d95dd3", 
    x"39d946c3", 
    x"39d92fb9", 
    x"39d918b3", 
    x"39d901b2", 
    x"39d8eab6", 
    x"39d8d3bf", 
    x"39d8bccc", 
    x"39d8a5df", 
    x"39d88ef6", 
    x"39d87813", 
    x"39d86134", 
    x"39d84a5a", 
    x"39d83384", 
    x"39d81cb4", 
    x"39d805e8", 
    x"39d7ef21", 
    x"39d7d85f", 
    x"39d7c1a2", 
    x"39d7aaea", 
    x"39d79436", 
    x"39d77d87", 
    x"39d766dd", 
    x"39d75038", 
    x"39d73997", 
    x"39d722fb", 
    x"39d70c64", 
    x"39d6f5d2", 
    x"39d6df44", 
    x"39d6c8bb", 
    x"39d6b237", 
    x"39d69bb7", 
    x"39d6853d", 
    x"39d66ec7", 
    x"39d65855", 
    x"39d641e9", 
    x"39d62b81", 
    x"39d6151e", 
    x"39d5febf", 
    x"39d5e865", 
    x"39d5d210", 
    x"39d5bbbf", 
    x"39d5a573", 
    x"39d58f2c", 
    x"39d578e9", 
    x"39d562ac", 
    x"39d54c72", 
    x"39d5363d", 
    x"39d5200d", 
    x"39d509e2", 
    x"39d4f3bb", 
    x"39d4dd99", 
    x"39d4c77b", 
    x"39d4b162", 
    x"39d49b4d", 
    x"39d4853e", 
    x"39d46f32", 
    x"39d4592b", 
    x"39d44329", 
    x"39d42d2c", 
    x"39d41733", 
    x"39d4013e", 
    x"39d3eb4e", 
    x"39d3d563", 
    x"39d3bf7c", 
    x"39d3a999", 
    x"39d393bb", 
    x"39d37de2", 
    x"39d3680d", 
    x"39d3523d", 
    x"39d33c71", 
    x"39d326aa", 
    x"39d310e7", 
    x"39d2fb28", 
    x"39d2e56f", 
    x"39d2cfb9", 
    x"39d2ba08", 
    x"39d2a45c", 
    x"39d28eb4", 
    x"39d27910", 
    x"39d26371", 
    x"39d24dd6", 
    x"39d23840", 
    x"39d222ae", 
    x"39d20d21", 
    x"39d1f798", 
    x"39d1e213", 
    x"39d1cc93", 
    x"39d1b717", 
    x"39d1a1a0", 
    x"39d18c2d", 
    x"39d176be", 
    x"39d16154", 
    x"39d14bee", 
    x"39d1368d", 
    x"39d12130", 
    x"39d10bd7", 
    x"39d0f683", 
    x"39d0e133", 
    x"39d0cbe7", 
    x"39d0b6a0", 
    x"39d0a15d", 
    x"39d08c1e", 
    x"39d076e4", 
    x"39d061ae", 
    x"39d04c7c", 
    x"39d0374f", 
    x"39d02226", 
    x"39d00d01", 
    x"39cff7e0", 
    x"39cfe2c4", 
    x"39cfcdac", 
    x"39cfb899", 
    x"39cfa389", 
    x"39cf8e7e", 
    x"39cf7977", 
    x"39cf6475", 
    x"39cf4f76", 
    x"39cf3a7c", 
    x"39cf2586", 
    x"39cf1095", 
    x"39cefba7", 
    x"39cee6be", 
    x"39ced1d9", 
    x"39cebcf9", 
    x"39cea81c", 
    x"39ce9344", 
    x"39ce7e70", 
    x"39ce69a0", 
    x"39ce54d4", 
    x"39ce400d", 
    x"39ce2b4a", 
    x"39ce168a", 
    x"39ce01d0", 
    x"39cded19", 
    x"39cdd866", 
    x"39cdc3b8", 
    x"39cdaf0d", 
    x"39cd9a67", 
    x"39cd85c5", 
    x"39cd7127", 
    x"39cd5c8e", 
    x"39cd47f8", 
    x"39cd3367", 
    x"39cd1ed9", 
    x"39cd0a50", 
    x"39ccf5cb", 
    x"39cce14a"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
