LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE target_fpga_pkg IS
    constant C_TARGET_DEVICE        : STRING := "U55";
end target_fpga_pkg;
