-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom1 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom1; 
 
architecture behavioral of inv_rom1 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"3b000000", 
    x"3aff8040", 
    x"3aff00ff", 
    x"3afe823d", 
    x"3afe03f8", 
    x"3afd8631", 
    x"3afd08e5", 
    x"3afc8c16", 
    x"3afc0fc1", 
    x"3afb93e6", 
    x"3afb1885", 
    x"3afa9d9d", 
    x"3afa232d", 
    x"3af9a934", 
    x"3af92fb2", 
    x"3af8b6a6", 
    x"3af83e10", 
    x"3af7c5ee", 
    x"3af74e40", 
    x"3af6d705", 
    x"3af6603e", 
    x"3af5e9e8", 
    x"3af57404", 
    x"3af4fe91", 
    x"3af4898d", 
    x"3af414fa", 
    x"3af3a0d5", 
    x"3af32d1f", 
    x"3af2b9d6", 
    x"3af246fb", 
    x"3af1d48c", 
    x"3af16289", 
    x"3af0f0f1", 
    x"3af07fc4", 
    x"3af00f01", 
    x"3aef9ea8", 
    x"3aef2eb7", 
    x"3aeebf2f", 
    x"3aee500f", 
    x"3aede156", 
    x"3aed7304", 
    x"3aed0518", 
    x"3aec9791", 
    x"3aec2a70", 
    x"3aebbdb3", 
    x"3aeb515a", 
    x"3aeae564", 
    x"3aea79d1", 
    x"3aea0ea1", 
    x"3ae9a3d2", 
    x"3ae93965", 
    x"3ae8cf59", 
    x"3ae865ac", 
    x"3ae7fc60", 
    x"3ae79373", 
    x"3ae72ae4", 
    x"3ae6c2b4", 
    x"3ae65ae2", 
    x"3ae5f36d", 
    x"3ae58c54", 
    x"3ae52598", 
    x"3ae4bf38", 
    x"3ae45933", 
    x"3ae3f389", 
    x"3ae38e39", 
    x"3ae32943", 
    x"3ae2c4a7", 
    x"3ae26063", 
    x"3ae1fc78", 
    x"3ae198e5", 
    x"3ae135aa", 
    x"3ae0d2c6", 
    x"3ae07038", 
    x"3ae00e01", 
    x"3adfac1f", 
    x"3adf4a93", 
    x"3adee95c", 
    x"3ade887a", 
    x"3ade27eb", 
    x"3addc7b0", 
    x"3add67c9", 
    x"3add0834", 
    x"3adca8f1", 
    x"3adc4a01", 
    x"3adbeb62", 
    x"3adb8d14", 
    x"3adb2f17", 
    x"3adad16a", 
    x"3ada740e", 
    x"3ada1700", 
    x"3ad9ba42", 
    x"3ad95dd3", 
    x"3ad901b2", 
    x"3ad8a5df", 
    x"3ad84a5a", 
    x"3ad7ef21", 
    x"3ad79436", 
    x"3ad73997", 
    x"3ad6df44", 
    x"3ad6853d", 
    x"3ad62b81", 
    x"3ad5d210", 
    x"3ad578e9", 
    x"3ad5200d", 
    x"3ad4c77b", 
    x"3ad46f32", 
    x"3ad41733", 
    x"3ad3bf7c", 
    x"3ad3680d", 
    x"3ad310e7", 
    x"3ad2ba08", 
    x"3ad26371", 
    x"3ad20d21", 
    x"3ad1b717", 
    x"3ad16154", 
    x"3ad10bd7", 
    x"3ad0b6a0", 
    x"3ad061ae", 
    x"3ad00d01", 
    x"3acfb899", 
    x"3acf6475", 
    x"3acf1095", 
    x"3acebcf9", 
    x"3ace69a0", 
    x"3ace168a", 
    x"3acdc3b8", 
    x"3acd7127", 
    x"3acd1ed9", 
    x"3acccccd", 
    x"3acc7b02", 
    x"3acc2978", 
    x"3acbd830", 
    x"3acb8728", 
    x"3acb3660", 
    x"3acae5d8", 
    x"3aca9590", 
    x"3aca4588", 
    x"3ac9f5bf", 
    x"3ac9a634", 
    x"3ac956e8", 
    x"3ac907da", 
    x"3ac8b90b", 
    x"3ac86a79", 
    x"3ac81c24", 
    x"3ac7ce0c", 
    x"3ac78032", 
    x"3ac73294", 
    x"3ac6e532", 
    x"3ac6980c", 
    x"3ac64b22", 
    x"3ac5fe74", 
    x"3ac5b201", 
    x"3ac565c8", 
    x"3ac519cb", 
    x"3ac4ce08", 
    x"3ac4827f", 
    x"3ac43730", 
    x"3ac3ec1a", 
    x"3ac3a13e", 
    x"3ac3569b", 
    x"3ac30c31", 
    x"3ac2c1ff", 
    x"3ac27806", 
    x"3ac22e45", 
    x"3ac1e4bc", 
    x"3ac19b6a", 
    x"3ac15250", 
    x"3ac1096d", 
    x"3ac0c0c1", 
    x"3ac0784b", 
    x"3ac0300c", 
    x"3abfe803", 
    x"3abfa030", 
    x"3abf5892", 
    x"3abf112b", 
    x"3abec9f8", 
    x"3abe82fa", 
    x"3abe3c31", 
    x"3abdf59d", 
    x"3abdaf3c", 
    x"3abd6910", 
    x"3abd2318", 
    x"3abcdd53", 
    x"3abc97c2", 
    x"3abc5264", 
    x"3abc0d39", 
    x"3abbc841", 
    x"3abb837b", 
    x"3abb3ee7", 
    x"3abafa86", 
    x"3abab656", 
    x"3aba7258", 
    x"3aba2e8c", 
    x"3ab9eaf0", 
    x"3ab9a786", 
    x"3ab9644d", 
    x"3ab92144", 
    x"3ab8de6c", 
    x"3ab89bc3", 
    x"3ab8594b", 
    x"3ab81703", 
    x"3ab7d4ea", 
    x"3ab79301", 
    x"3ab75147", 
    x"3ab70fbb", 
    x"3ab6ce5f", 
    x"3ab68d31", 
    x"3ab64c32", 
    x"3ab60b61", 
    x"3ab5cabe", 
    x"3ab58a48", 
    x"3ab54a01", 
    x"3ab509e7", 
    x"3ab4c9fa", 
    x"3ab48a3a", 
    x"3ab44aa7", 
    x"3ab40b41", 
    x"3ab3cc07", 
    x"3ab38cfa", 
    x"3ab34e19", 
    x"3ab30f63", 
    x"3ab2d0da", 
    x"3ab2927c", 
    x"3ab2544a", 
    x"3ab21643", 
    x"3ab1d867", 
    x"3ab19ab6", 
    x"3ab15d2f", 
    x"3ab11fd4", 
    x"3ab0e2a2", 
    x"3ab0a59b", 
    x"3ab068be", 
    x"3ab02c0b", 
    x"3aafef82", 
    x"3aafb322", 
    x"3aaf76eb", 
    x"3aaf3ade", 
    x"3aaefefa", 
    x"3aaec33e", 
    x"3aae87ab", 
    x"3aae4c41", 
    x"3aae1100", 
    x"3aadd5e6", 
    x"3aad9af5", 
    x"3aad602b", 
    x"3aad258a", 
    x"3aaceb10", 
    x"3aacb0bd", 
    x"3aac7692", 
    x"3aac3c8d", 
    x"3aac02b0", 
    x"3aabc8fa", 
    x"3aab8f6a", 
    x"3aab5601", 
    x"3aab1cbe", 
    x"3aaae3a1", 
    x"3aaaaaab", 
    x"3aaa71da", 
    x"3aaa392f", 
    x"3aaa00aa", 
    x"3aa9c84a", 
    x"3aa99010", 
    x"3aa957fb", 
    x"3aa9200b", 
    x"3aa8e83f", 
    x"3aa8b099", 
    x"3aa87917", 
    x"3aa841ba", 
    x"3aa80a81", 
    x"3aa7d36c", 
    x"3aa79c7b", 
    x"3aa765ae", 
    x"3aa72f05", 
    x"3aa6f880", 
    x"3aa6c21e", 
    x"3aa68bdf", 
    x"3aa655c4", 
    x"3aa61fcc", 
    x"3aa5e9f7", 
    x"3aa5b445", 
    x"3aa57eb5", 
    x"3aa54948", 
    x"3aa513fd", 
    x"3aa4ded5", 
    x"3aa4a9cf", 
    x"3aa474eb", 
    x"3aa44029", 
    x"3aa40b89", 
    x"3aa3d70a", 
    x"3aa3a2ad", 
    x"3aa36e72", 
    x"3aa33a57", 
    x"3aa3065e", 
    x"3aa2d286", 
    x"3aa29ecf", 
    x"3aa26b39", 
    x"3aa237c3", 
    x"3aa2046e", 
    x"3aa1d13a", 
    x"3aa19e25", 
    x"3aa16b31", 
    x"3aa1385d", 
    x"3aa105a9", 
    x"3aa0d315", 
    x"3aa0a0a1", 
    x"3aa06e4c", 
    x"3aa03c17", 
    x"3aa00a01", 
    x"3a9fd80a", 
    x"3a9fa633", 
    x"3a9f747a", 
    x"3a9f42e1", 
    x"3a9f1166", 
    x"3a9ee00a", 
    x"3a9eaecd", 
    x"3a9e7dae", 
    x"3a9e4cad", 
    x"3a9e1bcb", 
    x"3a9deb07", 
    x"3a9dba61", 
    x"3a9d89d9", 
    x"3a9d596e", 
    x"3a9d2922", 
    x"3a9cf8f3", 
    x"3a9cc8e1", 
    x"3a9c98ed", 
    x"3a9c6917", 
    x"3a9c395d", 
    x"3a9c09c1", 
    x"3a9bda41", 
    x"3a9baadf", 
    x"3a9b7b99", 
    x"3a9b4c70", 
    x"3a9b1d63", 
    x"3a9aee73", 
    x"3a9abf9f", 
    x"3a9a90e8", 
    x"3a9a624d", 
    x"3a9a33cd", 
    x"3a9a056a", 
    x"3a99d723", 
    x"3a99a8f7", 
    x"3a997ae7", 
    x"3a994cf3", 
    x"3a991f1a", 
    x"3a98f15d", 
    x"3a98c3bb", 
    x"3a989634", 
    x"3a9868c8", 
    x"3a983b77", 
    x"3a980e41", 
    x"3a97e126", 
    x"3a97b426", 
    x"3a978740", 
    x"3a975a75", 
    x"3a972dc4", 
    x"3a97012e", 
    x"3a96d4b2", 
    x"3a96a850", 
    x"3a967c08", 
    x"3a964fda", 
    x"3a9623c7", 
    x"3a95f7cc", 
    x"3a95cbec", 
    x"3a95a025", 
    x"3a957478", 
    x"3a9548e5", 
    x"3a951d6a", 
    x"3a94f209", 
    x"3a94c6c2", 
    x"3a949b93", 
    x"3a94707d", 
    x"3a944581", 
    x"3a941a9d", 
    x"3a93efd2", 
    x"3a93c51f", 
    x"3a939a86", 
    x"3a937005", 
    x"3a93459c", 
    x"3a931b4c", 
    x"3a92f114", 
    x"3a92c6f4", 
    x"3a929cec", 
    x"3a9272fc", 
    x"3a924925", 
    x"3a921f65", 
    x"3a91f5bd", 
    x"3a91cc2c", 
    x"3a91a2b4", 
    x"3a917953", 
    x"3a915009", 
    x"3a9126d7", 
    x"3a90fdbc", 
    x"3a90d4b8", 
    x"3a90abcc", 
    x"3a9082f7", 
    x"3a905a38", 
    x"3a903191", 
    x"3a900901", 
    x"3a8fe087", 
    x"3a8fb824", 
    x"3a8f8fd8", 
    x"3a8f67a2", 
    x"3a8f3f83", 
    x"3a8f177a", 
    x"3a8eef87", 
    x"3a8ec7ab", 
    x"3a8e9fe5", 
    x"3a8e7835", 
    x"3a8e509c", 
    x"3a8e2918", 
    x"3a8e01aa", 
    x"3a8dda52", 
    x"3a8db310", 
    x"3a8d8be3", 
    x"3a8d64cc", 
    x"3a8d3dcb", 
    x"3a8d16df", 
    x"3a8cf009", 
    x"3a8cc948", 
    x"3a8ca29c", 
    x"3a8c7c05", 
    x"3a8c5584", 
    x"3a8c2f18", 
    x"3a8c08c1", 
    x"3a8be27e", 
    x"3a8bbc51", 
    x"3a8b9638", 
    x"3a8b7034", 
    x"3a8b4a45", 
    x"3a8b246b", 
    x"3a8afea5", 
    x"3a8ad8f3", 
    x"3a8ab356", 
    x"3a8a8dcd", 
    x"3a8a6859", 
    x"3a8a42f8", 
    x"3a8a1dac", 
    x"3a89f874", 
    x"3a89d350", 
    x"3a89ae41", 
    x"3a898944", 
    x"3a89645c", 
    x"3a893f88", 
    x"3a891ac7", 
    x"3a88f61a", 
    x"3a88d181", 
    x"3a88acfb", 
    x"3a888889", 
    x"3a88642a", 
    x"3a883fde", 
    x"3a881ba6", 
    x"3a87f781", 
    x"3a87d36f", 
    x"3a87af70", 
    x"3a878b84", 
    x"3a8767ab", 
    x"3a8743e6", 
    x"3a872033", 
    x"3a86fc93", 
    x"3a86d905", 
    x"3a86b58b", 
    x"3a869223", 
    x"3a866ecd", 
    x"3a864b8a", 
    x"3a86285a", 
    x"3a86053c", 
    x"3a85e231", 
    x"3a85bf37", 
    x"3a859c50", 
    x"3a85797c", 
    x"3a8556b9", 
    x"3a853408", 
    x"3a85116a", 
    x"3a84eedd", 
    x"3a84cc63", 
    x"3a84a9fa", 
    x"3a8487a3", 
    x"3a84655e", 
    x"3a84432a", 
    x"3a842108", 
    x"3a83fef8", 
    x"3a83dcf9", 
    x"3a83bb0c", 
    x"3a839930", 
    x"3a837766", 
    x"3a8355ad", 
    x"3a833405", 
    x"3a83126f", 
    x"3a82f0e9", 
    x"3a82cf75", 
    x"3a82ae12", 
    x"3a828cc0", 
    x"3a826b7f", 
    x"3a824a4e", 
    x"3a82292f", 
    x"3a820821", 
    x"3a81e723", 
    x"3a81c636", 
    x"3a81a559", 
    x"3a81848e", 
    x"3a8163d3", 
    x"3a814328", 
    x"3a81228e", 
    x"3a810204", 
    x"3a80e18b", 
    x"3a80c122", 
    x"3a80a0c9", 
    x"3a808081", 
    x"3a806048", 
    x"3a804020", 
    x"3a802008"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
