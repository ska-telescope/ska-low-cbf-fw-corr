-- Created by python script create_inv_roms.py 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity inv_rom7 is 
port( 
    i_clk  : in  std_logic; 
    i_addr : in  std_logic_vector(8 downto 0); 
    o_data : out std_logic_vector(31 downto 0) 
    ); 
end inv_rom7; 
 
architecture behavioral of inv_rom7 is 
    type rom_type is array(511 downto 0) of std_logic_vector(31 downto 0); 
    signal rom : rom_type := (
    x"39800801", 
    x"39801002", 
    x"39801805", 
    x"39802008", 
    x"3980280d", 
    x"39803012", 
    x"39803819", 
    x"39804020", 
    x"39804829", 
    x"39805032", 
    x"3980583d", 
    x"39806048", 
    x"39806855", 
    x"39807062", 
    x"39807871", 
    x"39808081", 
    x"39808891", 
    x"398090a3", 
    x"398098b5", 
    x"3980a0c9", 
    x"3980a8de", 
    x"3980b0f3", 
    x"3980b90a", 
    x"3980c122", 
    x"3980c93a", 
    x"3980d154", 
    x"3980d96f", 
    x"3980e18b", 
    x"3980e9a7", 
    x"3980f1c5", 
    x"3980f9e4", 
    x"39810204", 
    x"39810a25", 
    x"39811247", 
    x"39811a6a", 
    x"3981228e", 
    x"39812ab3", 
    x"398132d9", 
    x"39813b00", 
    x"39814328", 
    x"39814b51", 
    x"3981537b", 
    x"39815ba6", 
    x"398163d3", 
    x"39816c00", 
    x"3981742e", 
    x"39817c5d", 
    x"3981848e", 
    x"39818cbf", 
    x"398194f1", 
    x"39819d25", 
    x"3981a559", 
    x"3981ad8f", 
    x"3981b5c5", 
    x"3981bdfd", 
    x"3981c636", 
    x"3981ce6f", 
    x"3981d6aa", 
    x"3981dee6", 
    x"3981e723", 
    x"3981ef61", 
    x"3981f7a0", 
    x"3981ffe0", 
    x"39820821", 
    x"39821063", 
    x"398218a6", 
    x"398220ea", 
    x"3982292f", 
    x"39823175", 
    x"398239bd", 
    x"39824205", 
    x"39824a4e", 
    x"39825299", 
    x"39825ae4", 
    x"39826331", 
    x"39826b7f", 
    x"398273cd", 
    x"39827c1d", 
    x"3982846e", 
    x"39828cc0", 
    x"39829513", 
    x"39829d67", 
    x"3982a5bc", 
    x"3982ae12", 
    x"3982b669", 
    x"3982bec1", 
    x"3982c71b", 
    x"3982cf75", 
    x"3982d7d0", 
    x"3982e02d", 
    x"3982e88b", 
    x"3982f0e9", 
    x"3982f949", 
    x"398301aa", 
    x"39830a0c", 
    x"3983126f", 
    x"39831ad3", 
    x"39832338", 
    x"39832b9e", 
    x"39833405", 
    x"39833c6d", 
    x"398344d7", 
    x"39834d41", 
    x"398355ad", 
    x"39835e1a", 
    x"39836687", 
    x"39836ef6", 
    x"39837766", 
    x"39837fd7", 
    x"39838849", 
    x"398390bc", 
    x"39839930", 
    x"3983a1a6", 
    x"3983aa1c", 
    x"3983b294", 
    x"3983bb0c", 
    x"3983c386", 
    x"3983cc01", 
    x"3983d47c", 
    x"3983dcf9", 
    x"3983e577", 
    x"3983edf6", 
    x"3983f677", 
    x"3983fef8", 
    x"3984077a", 
    x"39840ffe", 
    x"39841883", 
    x"39842108", 
    x"3984298f", 
    x"39843217", 
    x"39843aa0", 
    x"3984432a", 
    x"39844bb5", 
    x"39845442", 
    x"39845ccf", 
    x"3984655e", 
    x"39846ded", 
    x"3984767e", 
    x"39847f10", 
    x"398487a3", 
    x"39849037", 
    x"398498cc", 
    x"3984a162", 
    x"3984a9fa", 
    x"3984b292", 
    x"3984bb2c", 
    x"3984c3c7", 
    x"3984cc63", 
    x"3984d500", 
    x"3984dd9e", 
    x"3984e63d", 
    x"3984eedd", 
    x"3984f77f", 
    x"39850021", 
    x"398508c5", 
    x"3985116a", 
    x"39851a10", 
    x"398522b7", 
    x"39852b5f", 
    x"39853408", 
    x"39853cb3", 
    x"3985455e", 
    x"39854e0b", 
    x"398556b9", 
    x"39855f68", 
    x"39856818", 
    x"398570c9", 
    x"3985797c", 
    x"3985822f", 
    x"39858ae4", 
    x"39859399", 
    x"39859c50", 
    x"3985a508", 
    x"3985adc2", 
    x"3985b67c", 
    x"3985bf37", 
    x"3985c7f4", 
    x"3985d0b2", 
    x"3985d971", 
    x"3985e231", 
    x"3985eaf2", 
    x"3985f3b4", 
    x"3985fc78", 
    x"3986053c", 
    x"39860e02", 
    x"398616c9", 
    x"39861f91", 
    x"3986285a", 
    x"39863124", 
    x"398639f0", 
    x"398642bd", 
    x"39864b8a", 
    x"39865459", 
    x"39865d2a", 
    x"398665fb", 
    x"39866ecd", 
    x"398677a1", 
    x"39868076", 
    x"3986894c", 
    x"39869223", 
    x"39869afb", 
    x"3986a3d4", 
    x"3986acaf", 
    x"3986b58b", 
    x"3986be68", 
    x"3986c746", 
    x"3986d025", 
    x"3986d905", 
    x"3986e1e7", 
    x"3986eaca", 
    x"3986f3ae", 
    x"3986fc93", 
    x"39870579", 
    x"39870e60", 
    x"39871749", 
    x"39872033", 
    x"3987291e", 
    x"3987320a", 
    x"39873af7", 
    x"398743e6", 
    x"39874cd5", 
    x"398755c6", 
    x"39875eb8", 
    x"398767ab", 
    x"398770a0", 
    x"39877995", 
    x"3987828c", 
    x"39878b84", 
    x"3987947d", 
    x"39879d78", 
    x"3987a673", 
    x"3987af70", 
    x"3987b86e", 
    x"3987c16d", 
    x"3987ca6d", 
    x"3987d36f", 
    x"3987dc71", 
    x"3987e575", 
    x"3987ee7a", 
    x"3987f781", 
    x"39880088", 
    x"39880991", 
    x"3988129b", 
    x"39881ba6", 
    x"398824b2", 
    x"39882dbf", 
    x"398836ce", 
    x"39883fde", 
    x"398848ef", 
    x"39885201", 
    x"39885b15", 
    x"3988642a", 
    x"39886d3f", 
    x"39887657", 
    x"39887f6f", 
    x"39888889", 
    x"398891a3", 
    x"39889abf", 
    x"3988a3dd", 
    x"3988acfb", 
    x"3988b61b", 
    x"3988bf3b", 
    x"3988c85e", 
    x"3988d181", 
    x"3988daa5", 
    x"3988e3cb", 
    x"3988ecf2", 
    x"3988f61a", 
    x"3988ff44", 
    x"3989086e", 
    x"3989119a", 
    x"39891ac7", 
    x"398923f6", 
    x"39892d25", 
    x"39893656", 
    x"39893f88", 
    x"398948bb", 
    x"398951f0", 
    x"39895b25", 
    x"3989645c", 
    x"39896d95", 
    x"398976ce", 
    x"39898009", 
    x"39898944", 
    x"39899282", 
    x"39899bc0", 
    x"3989a500", 
    x"3989ae41", 
    x"3989b783", 
    x"3989c0c6", 
    x"3989ca0b", 
    x"3989d350", 
    x"3989dc98", 
    x"3989e5e0", 
    x"3989ef2a", 
    x"3989f874", 
    x"398a01c1", 
    x"398a0b0e", 
    x"398a145d", 
    x"398a1dac", 
    x"398a26fe", 
    x"398a3050", 
    x"398a39a4", 
    x"398a42f8", 
    x"398a4c4f", 
    x"398a55a6", 
    x"398a5eff", 
    x"398a6859", 
    x"398a71b4", 
    x"398a7b10", 
    x"398a846e", 
    x"398a8dcd", 
    x"398a972d", 
    x"398aa08f", 
    x"398aa9f2", 
    x"398ab356", 
    x"398abcbb", 
    x"398ac622", 
    x"398acf8a", 
    x"398ad8f3", 
    x"398ae25d", 
    x"398aebc9", 
    x"398af536", 
    x"398afea5", 
    x"398b0814", 
    x"398b1185", 
    x"398b1af7", 
    x"398b246b", 
    x"398b2ddf", 
    x"398b3755", 
    x"398b40cd", 
    x"398b4a45", 
    x"398b53bf", 
    x"398b5d3a", 
    x"398b66b7", 
    x"398b7034", 
    x"398b79b3", 
    x"398b8334", 
    x"398b8cb5", 
    x"398b9638", 
    x"398b9fbc", 
    x"398ba942", 
    x"398bb2c9", 
    x"398bbc51", 
    x"398bc5da", 
    x"398bcf65", 
    x"398bd8f1", 
    x"398be27e", 
    x"398bec0d", 
    x"398bf59d", 
    x"398bff2e", 
    x"398c08c1", 
    x"398c1254", 
    x"398c1bea", 
    x"398c2580", 
    x"398c2f18", 
    x"398c38b1", 
    x"398c424b", 
    x"398c4be7", 
    x"398c5584", 
    x"398c5f22", 
    x"398c68c2", 
    x"398c7263", 
    x"398c7c05", 
    x"398c85a9", 
    x"398c8f4e", 
    x"398c98f4", 
    x"398ca29c", 
    x"398cac45", 
    x"398cb5ef", 
    x"398cbf9b", 
    x"398cc948", 
    x"398cd2f6", 
    x"398cdca6", 
    x"398ce657", 
    x"398cf009", 
    x"398cf9bc", 
    x"398d0371", 
    x"398d0d28", 
    x"398d16df", 
    x"398d2098", 
    x"398d2a52", 
    x"398d340e", 
    x"398d3dcb", 
    x"398d4789", 
    x"398d5149", 
    x"398d5b0a", 
    x"398d64cc", 
    x"398d6e90", 
    x"398d7855", 
    x"398d821c", 
    x"398d8be3", 
    x"398d95ac", 
    x"398d9f77", 
    x"398da943", 
    x"398db310", 
    x"398dbcde", 
    x"398dc6ae", 
    x"398dd07f", 
    x"398dda52", 
    x"398de426", 
    x"398dedfb", 
    x"398df7d2", 
    x"398e01aa", 
    x"398e0b83", 
    x"398e155e", 
    x"398e1f3a", 
    x"398e2918", 
    x"398e32f7", 
    x"398e3cd7", 
    x"398e46b9", 
    x"398e509c", 
    x"398e5a80", 
    x"398e6466", 
    x"398e6e4d", 
    x"398e7835", 
    x"398e821f", 
    x"398e8c0b", 
    x"398e95f7", 
    x"398e9fe5", 
    x"398ea9d5", 
    x"398eb3c5", 
    x"398ebdb8", 
    x"398ec7ab", 
    x"398ed1a0", 
    x"398edb97", 
    x"398ee58e", 
    x"398eef87", 
    x"398ef982", 
    x"398f037e", 
    x"398f0d7b", 
    x"398f177a", 
    x"398f217a", 
    x"398f2b7b", 
    x"398f357e", 
    x"398f3f83", 
    x"398f4988", 
    x"398f538f", 
    x"398f5d98", 
    x"398f67a2", 
    x"398f71ad", 
    x"398f7bba", 
    x"398f85c8", 
    x"398f8fd8", 
    x"398f99e9", 
    x"398fa3fb", 
    x"398fae0f", 
    x"398fb824", 
    x"398fc23b", 
    x"398fcc53", 
    x"398fd66c", 
    x"398fe087", 
    x"398feaa3", 
    x"398ff4c1", 
    x"398ffee0", 
    x"39900901", 
    x"39901323", 
    x"39901d46", 
    x"3990276b", 
    x"39903191", 
    x"39903bb9", 
    x"399045e2", 
    x"3990500c", 
    x"39905a38", 
    x"39906466", 
    x"39906e95", 
    x"399078c5", 
    x"399082f7", 
    x"39908d2a", 
    x"3990975e", 
    x"3990a195", 
    x"3990abcc", 
    x"3990b605", 
    x"3990c03f", 
    x"3990ca7b", 
    x"3990d4b8", 
    x"3990def7", 
    x"3990e937", 
    x"3990f379", 
    x"3990fdbc", 
    x"39910801", 
    x"39911247", 
    x"39911c8e", 
    x"399126d7", 
    x"39913121", 
    x"39913b6d", 
    x"399145ba", 
    x"39915009", 
    x"39915a59", 
    x"399164ab", 
    x"39916efe", 
    x"39917953", 
    x"399183a9", 
    x"39918e00", 
    x"39919859", 
    x"3991a2b4", 
    x"3991ad10", 
    x"3991b76d", 
    x"3991c1cc", 
    x"3991cc2c", 
    x"3991d68e", 
    x"3991e0f2", 
    x"3991eb56", 
    x"3991f5bd", 
    x"39920025", 
    x"39920a8e", 
    x"399214f9", 
    x"39921f65", 
    x"399229d2", 
    x"39923442", 
    x"39923eb2", 
    x"39924925"); 
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
    signal data : std_logic_vector(31 downto 0);
    
begin 
    process(i_clk) 
    begin 
        if rising_edge(i_clk) then 
            data <= ROM(conv_integer(i_addr)); 
            o_data <= data;
        end if;
    end process;
end behavioral; 
